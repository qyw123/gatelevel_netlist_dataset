
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386;

  GTECH_MUX2 U140 ( .A(n279), .B(n280), .S(n281), .Z(sum[9]) );
  GTECH_XNOR2 U141 ( .A(n282), .B(n283), .Z(n280) );
  GTECH_XOR2 U142 ( .A(n282), .B(n284), .Z(n279) );
  GTECH_AOI21 U143 ( .A(a[9]), .B(b[9]), .C(n285), .Z(n282) );
  GTECH_NAND2 U144 ( .A(n286), .B(n287), .Z(sum[8]) );
  GTECH_OAI21 U145 ( .A(n284), .B(n283), .C(n281), .Z(n286) );
  GTECH_MUX2 U146 ( .A(n288), .B(n289), .S(n290), .Z(sum[7]) );
  GTECH_XNOR2 U147 ( .A(n291), .B(n292), .Z(n289) );
  GTECH_OA21 U148 ( .A(n293), .B(n294), .C(n295), .Z(n292) );
  GTECH_NOR2 U149 ( .A(b[6]), .B(a[6]), .Z(n293) );
  GTECH_XOR2 U150 ( .A(n291), .B(n296), .Z(n288) );
  GTECH_XOR2 U151 ( .A(a[7]), .B(b[7]), .Z(n291) );
  GTECH_OAI21 U152 ( .A(n297), .B(n295), .C(n298), .Z(sum[6]) );
  GTECH_MUX2 U153 ( .A(n299), .B(n300), .S(b[6]), .Z(n298) );
  GTECH_OR_NOT U154 ( .A(a[6]), .B(n297), .Z(n300) );
  GTECH_XOR2 U155 ( .A(a[6]), .B(n297), .Z(n299) );
  GTECH_OA21 U156 ( .A(n290), .B(n301), .C(n294), .Z(n297) );
  GTECH_AO21 U157 ( .A(n302), .B(n303), .C(n304), .Z(n294) );
  GTECH_XOR2 U158 ( .A(n305), .B(n306), .Z(sum[5]) );
  GTECH_AOI21 U159 ( .A(n302), .B(n290), .C(n307), .Z(n306) );
  GTECH_AND_NOT U160 ( .A(n303), .B(n304), .Z(n305) );
  GTECH_XOR2 U161 ( .A(n308), .B(n290), .Z(sum[4]) );
  GTECH_MUX2 U162 ( .A(n309), .B(n310), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U163 ( .A(n311), .B(n312), .Z(n310) );
  GTECH_XNOR2 U164 ( .A(n311), .B(n313), .Z(n309) );
  GTECH_OA21 U165 ( .A(n314), .B(n315), .C(n316), .Z(n313) );
  GTECH_NOR2 U166 ( .A(a[2]), .B(b[2]), .Z(n314) );
  GTECH_XOR2 U167 ( .A(a[3]), .B(b[3]), .Z(n311) );
  GTECH_MUX2 U168 ( .A(n317), .B(n318), .S(cin), .Z(sum[2]) );
  GTECH_MUX2 U169 ( .A(n319), .B(n320), .S(n321), .Z(n318) );
  GTECH_MUX2 U170 ( .A(n320), .B(n319), .S(n315), .Z(n317) );
  GTECH_OAI21 U171 ( .A(n322), .B(n323), .C(n324), .Z(n315) );
  GTECH_XOR2 U172 ( .A(a[2]), .B(b[2]), .Z(n319) );
  GTECH_OAI21 U173 ( .A(b[2]), .B(a[2]), .C(n316), .Z(n320) );
  GTECH_MUX2 U174 ( .A(n325), .B(n326), .S(n327), .Z(sum[1]) );
  GTECH_AND_NOT U175 ( .A(n324), .B(n322), .Z(n327) );
  GTECH_OAI21 U176 ( .A(cin), .B(n323), .C(n328), .Z(n326) );
  GTECH_AO21 U177 ( .A(n328), .B(cin), .C(n323), .Z(n325) );
  GTECH_ADD_AB U178 ( .A(a[0]), .B(b[0]), .COUT(n323) );
  GTECH_MUX2 U179 ( .A(n329), .B(n330), .S(n331), .Z(sum[15]) );
  GTECH_XOR2 U180 ( .A(n332), .B(n333), .Z(n330) );
  GTECH_OA21 U181 ( .A(n334), .B(n335), .C(n336), .Z(n333) );
  GTECH_AND_NOT U182 ( .A(n337), .B(n338), .Z(n334) );
  GTECH_XNOR2 U183 ( .A(n332), .B(n339), .Z(n329) );
  GTECH_XNOR2 U184 ( .A(a[15]), .B(b[15]), .Z(n332) );
  GTECH_OAI21 U185 ( .A(n340), .B(n336), .C(n341), .Z(sum[14]) );
  GTECH_MUX2 U186 ( .A(n342), .B(n343), .S(b[14]), .Z(n341) );
  GTECH_OR_NOT U187 ( .A(a[14]), .B(n340), .Z(n343) );
  GTECH_XOR2 U188 ( .A(a[14]), .B(n340), .Z(n342) );
  GTECH_OA21 U189 ( .A(n344), .B(n345), .C(n337), .Z(n340) );
  GTECH_AOI21 U190 ( .A(n346), .B(n347), .C(n338), .Z(n345) );
  GTECH_MUX2 U191 ( .A(n348), .B(n349), .S(n331), .Z(sum[13]) );
  GTECH_XNOR2 U192 ( .A(n350), .B(n351), .Z(n349) );
  GTECH_XNOR2 U193 ( .A(n352), .B(n350), .Z(n348) );
  GTECH_AND_NOT U194 ( .A(n337), .B(n344), .Z(n350) );
  GTECH_NOT U195 ( .A(n353), .Z(n344) );
  GTECH_NAND2 U196 ( .A(n354), .B(n355), .Z(sum[12]) );
  GTECH_AO21 U197 ( .A(n351), .B(n347), .C(n331), .Z(n354) );
  GTECH_NOT U198 ( .A(n352), .Z(n347) );
  GTECH_NOT U199 ( .A(n338), .Z(n351) );
  GTECH_MUX2 U200 ( .A(n356), .B(n357), .S(n281), .Z(sum[11]) );
  GTECH_XOR2 U201 ( .A(n358), .B(n359), .Z(n357) );
  GTECH_XNOR2 U202 ( .A(n358), .B(n360), .Z(n356) );
  GTECH_OA21 U203 ( .A(n361), .B(n362), .C(n363), .Z(n360) );
  GTECH_ADD_AB U204 ( .A(n364), .B(n365), .COUT(n361) );
  GTECH_XOR2 U205 ( .A(a[11]), .B(b[11]), .Z(n358) );
  GTECH_OAI21 U206 ( .A(n366), .B(n363), .C(n367), .Z(sum[10]) );
  GTECH_MUX2 U207 ( .A(n368), .B(n369), .S(b[10]), .Z(n367) );
  GTECH_NAND2 U208 ( .A(n365), .B(n366), .Z(n369) );
  GTECH_XOR2 U209 ( .A(a[10]), .B(n366), .Z(n368) );
  GTECH_OA21 U210 ( .A(n370), .B(n371), .C(n362), .Z(n366) );
  GTECH_AOI2N2 U211 ( .A(a[9]), .B(b[9]), .C(n285), .D(n372), .Z(n362) );
  GTECH_NOT U212 ( .A(n284), .Z(n372) );
  GTECH_XNOR2 U213 ( .A(cin), .B(n373), .Z(sum[0]) );
  GTECH_OAI21 U214 ( .A(n331), .B(n374), .C(n355), .Z(cout) );
  GTECH_OR3 U215 ( .A(n338), .B(n352), .C(n346), .Z(n355) );
  GTECH_ADD_AB U216 ( .A(a[12]), .B(b[12]), .COUT(n338) );
  GTECH_AOI21 U217 ( .A(n339), .B(a[15]), .C(n375), .Z(n374) );
  GTECH_OA21 U218 ( .A(a[15]), .B(n339), .C(b[15]), .Z(n375) );
  GTECH_NAND2 U219 ( .A(n376), .B(n336), .Z(n339) );
  GTECH_NAND2 U220 ( .A(b[14]), .B(a[14]), .Z(n336) );
  GTECH_AO21 U221 ( .A(n337), .B(n352), .C(n335), .Z(n376) );
  GTECH_OAI21 U222 ( .A(b[14]), .B(a[14]), .C(n353), .Z(n335) );
  GTECH_OR2 U223 ( .A(b[13]), .B(a[13]), .Z(n353) );
  GTECH_NOR2 U224 ( .A(b[12]), .B(a[12]), .Z(n352) );
  GTECH_NAND2 U225 ( .A(a[13]), .B(b[13]), .Z(n337) );
  GTECH_NOT U226 ( .A(n346), .Z(n331) );
  GTECH_OAI21 U227 ( .A(n377), .B(n371), .C(n287), .Z(n346) );
  GTECH_OR3 U228 ( .A(n284), .B(n283), .C(n281), .Z(n287) );
  GTECH_NOT U229 ( .A(n371), .Z(n281) );
  GTECH_ADD_AB U230 ( .A(b[8]), .B(a[8]), .COUT(n284) );
  GTECH_MUX2 U231 ( .A(n378), .B(n308), .S(n290), .Z(n371) );
  GTECH_MUX2 U232 ( .A(n373), .B(n379), .S(cin), .Z(n290) );
  GTECH_AOI21 U233 ( .A(n312), .B(a[3]), .C(n380), .Z(n379) );
  GTECH_OA21 U234 ( .A(a[3]), .B(n312), .C(b[3]), .Z(n380) );
  GTECH_NAND2 U235 ( .A(n381), .B(n316), .Z(n312) );
  GTECH_NAND2 U236 ( .A(a[2]), .B(b[2]), .Z(n316) );
  GTECH_OAI21 U237 ( .A(a[2]), .B(b[2]), .C(n321), .Z(n381) );
  GTECH_OA21 U238 ( .A(n322), .B(n328), .C(n324), .Z(n321) );
  GTECH_OR2 U239 ( .A(a[1]), .B(b[1]), .Z(n324) );
  GTECH_OR2 U240 ( .A(a[0]), .B(b[0]), .Z(n328) );
  GTECH_ADD_AB U241 ( .A(b[1]), .B(a[1]), .COUT(n322) );
  GTECH_XNOR2 U242 ( .A(a[0]), .B(b[0]), .Z(n373) );
  GTECH_OR_NOT U243 ( .A(n307), .B(n302), .Z(n308) );
  GTECH_NAND2 U244 ( .A(b[4]), .B(a[4]), .Z(n302) );
  GTECH_AOI21 U245 ( .A(n296), .B(a[7]), .C(n382), .Z(n378) );
  GTECH_OA21 U246 ( .A(a[7]), .B(n296), .C(b[7]), .Z(n382) );
  GTECH_NAND2 U247 ( .A(n383), .B(n295), .Z(n296) );
  GTECH_NAND2 U248 ( .A(b[6]), .B(a[6]), .Z(n295) );
  GTECH_OAI21 U249 ( .A(a[6]), .B(b[6]), .C(n384), .Z(n383) );
  GTECH_NOT U250 ( .A(n301), .Z(n384) );
  GTECH_AO21 U251 ( .A(n303), .B(n307), .C(n304), .Z(n301) );
  GTECH_NOR2 U252 ( .A(a[5]), .B(b[5]), .Z(n304) );
  GTECH_NOR2 U253 ( .A(a[4]), .B(b[4]), .Z(n307) );
  GTECH_NAND2 U254 ( .A(b[5]), .B(a[5]), .Z(n303) );
  GTECH_AOI21 U255 ( .A(n359), .B(a[11]), .C(n385), .Z(n377) );
  GTECH_OA21 U256 ( .A(a[11]), .B(n359), .C(b[11]), .Z(n385) );
  GTECH_NAND2 U257 ( .A(n386), .B(n363), .Z(n359) );
  GTECH_OR_NOT U258 ( .A(n365), .B(b[10]), .Z(n363) );
  GTECH_AO21 U259 ( .A(n365), .B(n364), .C(n370), .Z(n386) );
  GTECH_AOI2N2 U260 ( .A(a[9]), .B(b[9]), .C(n283), .D(n285), .Z(n370) );
  GTECH_NOR2 U261 ( .A(b[9]), .B(a[9]), .Z(n285) );
  GTECH_NOR2 U262 ( .A(a[8]), .B(b[8]), .Z(n283) );
  GTECH_NOT U263 ( .A(b[10]), .Z(n364) );
  GTECH_NOT U264 ( .A(a[10]), .Z(n365) );
endmodule

