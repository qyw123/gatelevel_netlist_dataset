
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n111, n113, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n113), .K(n113), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n250) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n113), .K(n113), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n113), .K(n113), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n113), .K(n113), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n113), .K(n113), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n113), .K(n113), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]) );
  GTECH_FJK1S A_reg_15_ ( .J(n113), .K(n113), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n266) );
  GTECH_FJK1S A_reg_14_ ( .J(n113), .K(n113), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n265) );
  GTECH_FJK1S A_reg_13_ ( .J(n113), .K(n113), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n264) );
  GTECH_FJK1S A_reg_12_ ( .J(n113), .K(n113), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n263) );
  GTECH_FJK1S A_reg_11_ ( .J(n113), .K(n113), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n262) );
  GTECH_FJK1S A_reg_10_ ( .J(n113), .K(n113), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n261) );
  GTECH_FJK1S A_reg_9_ ( .J(n113), .K(n113), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n260) );
  GTECH_FJK1S A_reg_8_ ( .J(n113), .K(n113), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n259) );
  GTECH_FJK1S A_reg_7_ ( .J(n113), .K(n113), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n258) );
  GTECH_FJK1S A_reg_6_ ( .J(n113), .K(n113), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n257) );
  GTECH_FJK1S A_reg_5_ ( .J(n113), .K(n113), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n256) );
  GTECH_FJK1S A_reg_4_ ( .J(n113), .K(n113), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n255) );
  GTECH_FJK1S A_reg_3_ ( .J(n113), .K(n113), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n254) );
  GTECH_FJK1S A_reg_2_ ( .J(n113), .K(n113), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n253) );
  GTECH_FJK1S A_reg_1_ ( .J(n113), .K(n113), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n252) );
  GTECH_FJK1S A_reg_0_ ( .J(n113), .K(n113), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n251) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n113), .K(n113), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n113), .K(n113), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n113), .K(n113), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n113), .K(n113), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n113), .K(n113), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n113), .K(n113), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n113), .K(n113), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n113), .K(n113), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n113), .K(n113), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n113), .K(n113), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n113), .K(n113), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n113), .K(n113), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n113), .K(n113), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n113), .K(n113), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n113), .K(n113), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n113), .K(n113), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n113), .K(n113), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n113), .K(n113), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n113), .K(n113), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n113), .K(n113), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n113), .K(n113), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n113), .K(n113), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n113), .K(n113), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n113), .K(n113), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n113), .K(n113), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n113), .K(n113), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n113), .K(n113), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n113), .K(n113), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n113), .K(n113), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n113), .K(n113), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n113), .K(n113), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n113), .K(n113), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n113), .K(n113), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n113), .K(n113), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n113), .K(n113), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n113), .K(n113), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n113), .K(n113), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n113), .K(n113), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n113), .K(n113), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n113), .K(n113), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n113), .K(n113), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n113), .K(n113), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n113), .K(n113), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n113), .K(n113), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n113), .K(n113), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n113), .K(n113), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n113), .K(n113), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n113), .K(n113), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n113), .K(n113), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n113), .K(n113), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n113), .K(n113), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n113), .K(n113), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n113), .K(n113), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n113), .K(n113), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n113), .K(n113), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n113), .K(n113), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n113), .K(n113), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n113), .K(n113), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n113), .K(n113), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n113), .K(n113), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n113), .K(n113), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n113), .K(n113), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n113), .K(n113), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n113), .K(n113), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n113), .K(n113), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n113), .K(n113), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD2 Valid_reg ( .D(N155), .CP(clk), .CD(n111), .Q(Valid) );
  GTECH_ZERO U252 ( .Z(n113) );
  GTECH_ONE U253 ( .Z(n111) );
  GTECH_NOT U254 ( .A(n268), .Z(N99) );
  GTECH_AOI222 U255 ( .A(n269), .B(n270), .C(n271), .D(n272), .E(n273), .F(
        n274), .Z(n268) );
  GTECH_NOT U256 ( .A(n275), .Z(N98) );
  GTECH_AOI222 U257 ( .A(n271), .B(n276), .C(n277), .D(n278), .E(R[15]), .F(
        n279), .Z(n275) );
  GTECH_NAND2 U258 ( .A(n280), .B(n281), .Z(n277) );
  GTECH_OAI2N2 U259 ( .A(n13), .B(n282), .C(R[14]), .D(n279), .Z(N97) );
  GTECH_OAI2N2 U260 ( .A(n14), .B(n282), .C(R[13]), .D(n279), .Z(N96) );
  GTECH_OAI2N2 U261 ( .A(n15), .B(n282), .C(R[12]), .D(n279), .Z(N95) );
  GTECH_OAI2N2 U262 ( .A(n16), .B(n282), .C(R[11]), .D(n279), .Z(N94) );
  GTECH_OAI2N2 U263 ( .A(n17), .B(n282), .C(R[10]), .D(n279), .Z(N93) );
  GTECH_OAI2N2 U264 ( .A(n18), .B(n282), .C(R[9]), .D(n279), .Z(N92) );
  GTECH_OAI2N2 U265 ( .A(n19), .B(n282), .C(R[8]), .D(n279), .Z(N91) );
  GTECH_OAI2N2 U266 ( .A(n20), .B(n282), .C(R[7]), .D(n279), .Z(N90) );
  GTECH_OAI2N2 U267 ( .A(n21), .B(n282), .C(R[6]), .D(n279), .Z(N89) );
  GTECH_OAI2N2 U268 ( .A(n22), .B(n282), .C(R[5]), .D(n279), .Z(N88) );
  GTECH_OAI2N2 U269 ( .A(n23), .B(n282), .C(R[4]), .D(n279), .Z(N87) );
  GTECH_OAI2N2 U270 ( .A(n24), .B(n282), .C(R[3]), .D(n279), .Z(N86) );
  GTECH_OAI2N2 U271 ( .A(n25), .B(n282), .C(R[2]), .D(n279), .Z(N85) );
  GTECH_OAI2N2 U272 ( .A(n26), .B(n282), .C(R[1]), .D(n279), .Z(N84) );
  GTECH_OAI2N2 U273 ( .A(n27), .B(n282), .C(R[0]), .D(n279), .Z(N83) );
  GTECH_AND2 U274 ( .A(M[15]), .B(n279), .Z(N42) );
  GTECH_AND2 U275 ( .A(M[14]), .B(n279), .Z(N39) );
  GTECH_AND2 U276 ( .A(M[13]), .B(n279), .Z(N38) );
  GTECH_AND2 U277 ( .A(M[12]), .B(n279), .Z(N37) );
  GTECH_AND2 U278 ( .A(M[11]), .B(n279), .Z(N36) );
  GTECH_AND2 U279 ( .A(M[10]), .B(n279), .Z(N35) );
  GTECH_AND2 U280 ( .A(M[9]), .B(n279), .Z(N34) );
  GTECH_AND2 U281 ( .A(M[8]), .B(n279), .Z(N33) );
  GTECH_AND2 U282 ( .A(M[7]), .B(n279), .Z(N32) );
  GTECH_AND2 U283 ( .A(M[6]), .B(n279), .Z(N31) );
  GTECH_AND2 U284 ( .A(M[5]), .B(n279), .Z(N30) );
  GTECH_AND2 U285 ( .A(M[4]), .B(n279), .Z(N29) );
  GTECH_AND2 U286 ( .A(M[3]), .B(n279), .Z(N28) );
  GTECH_AND2 U287 ( .A(M[2]), .B(n279), .Z(N27) );
  GTECH_AND2 U288 ( .A(M[1]), .B(n279), .Z(N26) );
  GTECH_AND2 U289 ( .A(M[0]), .B(n279), .Z(N25) );
  GTECH_NOT U290 ( .A(n283), .Z(n279) );
  GTECH_NAND2 U291 ( .A(n283), .B(n284), .Z(N19) );
  GTECH_NAND3 U292 ( .A(n285), .B(n286), .C(n287), .Z(n284) );
  GTECH_NAND3 U293 ( .A(n288), .B(n289), .C(n282), .Z(N18) );
  GTECH_AND2 U294 ( .A(n287), .B(n290), .Z(N17) );
  GTECH_OAI21 U295 ( .A(n8), .B(n291), .C(n285), .Z(n290) );
  GTECH_AND2 U296 ( .A(n287), .B(n292), .Z(N16) );
  GTECH_OAI21 U297 ( .A(n7), .B(n293), .C(n294), .Z(n292) );
  GTECH_NOT U298 ( .A(n295), .Z(N152) );
  GTECH_AOI222 U299 ( .A(n296), .B(n297), .C(n298), .D(n299), .E(n300), .F(
        n301), .Z(n295) );
  GTECH_NAND2 U300 ( .A(n289), .B(n302), .Z(N151) );
  GTECH_NOT U301 ( .A(n303), .Z(N150) );
  GTECH_AOI222 U302 ( .A(n304), .B(n296), .C(n298), .D(n305), .E(n300), .F(
        n306), .Z(n303) );
  GTECH_MUX2 U303 ( .A(n307), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND_NOT U304 ( .A(n287), .B(n250), .Z(n307) );
  GTECH_NOT U305 ( .A(n308), .Z(N149) );
  GTECH_AOI222 U306 ( .A(n309), .B(n296), .C(n298), .D(n310), .E(n300), .F(
        n311), .Z(n308) );
  GTECH_NOT U307 ( .A(n312), .Z(N148) );
  GTECH_AOI222 U308 ( .A(n313), .B(n296), .C(n298), .D(n314), .E(n300), .F(
        n315), .Z(n312) );
  GTECH_NOT U309 ( .A(n316), .Z(N147) );
  GTECH_AOI222 U310 ( .A(n317), .B(n296), .C(n298), .D(n318), .E(n300), .F(
        n319), .Z(n316) );
  GTECH_NOT U311 ( .A(n320), .Z(N146) );
  GTECH_AOI222 U312 ( .A(n321), .B(n296), .C(n298), .D(n322), .E(n300), .F(
        n323), .Z(n320) );
  GTECH_NOT U313 ( .A(n324), .Z(N145) );
  GTECH_AOI222 U314 ( .A(n325), .B(n296), .C(n298), .D(n326), .E(n300), .F(
        n327), .Z(n324) );
  GTECH_NOT U315 ( .A(n328), .Z(N144) );
  GTECH_AOI222 U316 ( .A(n329), .B(n296), .C(n298), .D(n330), .E(n300), .F(
        n331), .Z(n328) );
  GTECH_NOT U317 ( .A(n332), .Z(N143) );
  GTECH_AOI222 U318 ( .A(n333), .B(n296), .C(n298), .D(n334), .E(n300), .F(
        n335), .Z(n332) );
  GTECH_NOT U319 ( .A(n336), .Z(N142) );
  GTECH_AOI222 U320 ( .A(n337), .B(n296), .C(n298), .D(n338), .E(n300), .F(
        n339), .Z(n336) );
  GTECH_NOT U321 ( .A(n340), .Z(N141) );
  GTECH_AOI222 U322 ( .A(n341), .B(n296), .C(n298), .D(n342), .E(n300), .F(
        n343), .Z(n340) );
  GTECH_NOT U323 ( .A(n344), .Z(N140) );
  GTECH_AOI222 U324 ( .A(n345), .B(n296), .C(n298), .D(n346), .E(n300), .F(
        n347), .Z(n344) );
  GTECH_NOT U325 ( .A(n348), .Z(N14) );
  GTECH_NAND2 U326 ( .A(n287), .B(n250), .Z(n348) );
  GTECH_NOT U327 ( .A(n349), .Z(N139) );
  GTECH_AOI222 U328 ( .A(n350), .B(n296), .C(n298), .D(n351), .E(n300), .F(
        n352), .Z(n349) );
  GTECH_NOT U329 ( .A(n353), .Z(N138) );
  GTECH_AOI222 U330 ( .A(n354), .B(n296), .C(n298), .D(n355), .E(n300), .F(
        n356), .Z(n353) );
  GTECH_NOT U331 ( .A(n357), .Z(N137) );
  GTECH_AOI222 U332 ( .A(n358), .B(n296), .C(n298), .D(n359), .E(n300), .F(
        n360), .Z(n357) );
  GTECH_NOT U333 ( .A(n361), .Z(N136) );
  GTECH_AOI222 U334 ( .A(n296), .B(n270), .C(n298), .D(n272), .E(n300), .F(
        n274), .Z(n361) );
  GTECH_NOT U335 ( .A(n362), .Z(n274) );
  GTECH_XOR2 U336 ( .A(n363), .B(n364), .Z(n362) );
  GTECH_NOT U337 ( .A(n365), .Z(n364) );
  GTECH_NOT U338 ( .A(n366), .Z(n298) );
  GTECH_NOT U339 ( .A(n367), .Z(n270) );
  GTECH_XOR2 U340 ( .A(n363), .B(n368), .Z(n367) );
  GTECH_NOT U341 ( .A(n369), .Z(n368) );
  GTECH_XOR2 U342 ( .A(n272), .B(n252), .Z(n363) );
  GTECH_OAI21 U343 ( .A(n12), .B(n366), .C(n370), .Z(N135) );
  GTECH_OAI21 U344 ( .A(n300), .B(n296), .C(n278), .Z(n370) );
  GTECH_OAI21 U345 ( .A(n12), .B(n371), .C(n365), .Z(n278) );
  GTECH_NOT U346 ( .A(n372), .Z(n296) );
  GTECH_NAND3 U347 ( .A(n28), .B(n373), .C(N155), .Z(n372) );
  GTECH_NOT U348 ( .A(n374), .Z(n300) );
  GTECH_NAND3 U349 ( .A(n10), .B(n375), .C(N155), .Z(n374) );
  GTECH_NAND2 U350 ( .A(n376), .B(N155), .Z(n366) );
  GTECH_XOR2 U351 ( .A(n373), .B(n28), .Z(n376) );
  GTECH_AND2 U352 ( .A(N155), .B(n377), .Z(N134) );
  GTECH_NOT U353 ( .A(n13), .Z(n377) );
  GTECH_AND2 U354 ( .A(N155), .B(n378), .Z(N133) );
  GTECH_NOT U355 ( .A(n14), .Z(n378) );
  GTECH_AND2 U356 ( .A(N155), .B(n379), .Z(N132) );
  GTECH_NOT U357 ( .A(n15), .Z(n379) );
  GTECH_AND2 U358 ( .A(N155), .B(n380), .Z(N131) );
  GTECH_NOT U359 ( .A(n16), .Z(n380) );
  GTECH_AND2 U360 ( .A(N155), .B(n381), .Z(N130) );
  GTECH_NOT U361 ( .A(n17), .Z(n381) );
  GTECH_AND2 U362 ( .A(N155), .B(n382), .Z(N129) );
  GTECH_NOT U363 ( .A(n18), .Z(n382) );
  GTECH_AND2 U364 ( .A(N155), .B(n383), .Z(N128) );
  GTECH_NOT U365 ( .A(n19), .Z(n383) );
  GTECH_AND2 U366 ( .A(N155), .B(n384), .Z(N127) );
  GTECH_NOT U367 ( .A(n20), .Z(n384) );
  GTECH_AND2 U368 ( .A(N155), .B(n385), .Z(N126) );
  GTECH_NOT U369 ( .A(n21), .Z(n385) );
  GTECH_AND2 U370 ( .A(N155), .B(n386), .Z(N125) );
  GTECH_NOT U371 ( .A(n22), .Z(n386) );
  GTECH_AND2 U372 ( .A(N155), .B(n387), .Z(N124) );
  GTECH_NOT U373 ( .A(n23), .Z(n387) );
  GTECH_AND2 U374 ( .A(N155), .B(n388), .Z(N123) );
  GTECH_NOT U375 ( .A(n24), .Z(n388) );
  GTECH_AND2 U376 ( .A(N155), .B(n389), .Z(N122) );
  GTECH_NOT U377 ( .A(n25), .Z(n389) );
  GTECH_AND2 U378 ( .A(N155), .B(n390), .Z(N121) );
  GTECH_NOT U379 ( .A(n26), .Z(n390) );
  GTECH_AND2 U380 ( .A(N155), .B(n391), .Z(N120) );
  GTECH_NOT U381 ( .A(n27), .Z(n391) );
  GTECH_NOT U382 ( .A(n302), .Z(N155) );
  GTECH_NAND5 U383 ( .A(n392), .B(n6), .C(n9), .D(n8), .E(n7), .Z(n302) );
  GTECH_NOR2 U384 ( .A(n250), .B(Rst), .Z(n392) );
  GTECH_NOT U385 ( .A(n393), .Z(N116) );
  GTECH_AOI222 U386 ( .A(n271), .B(n299), .C(n273), .D(n301), .E(n297), .F(
        n269), .Z(n393) );
  GTECH_XOR2 U387 ( .A(n394), .B(n395), .Z(n297) );
  GTECH_ADD_ABC U388 ( .A(n31), .B(n266), .C(n396), .COUT(n395) );
  GTECH_XOR2 U389 ( .A(n397), .B(n394), .Z(n301) );
  GTECH_XOR2 U390 ( .A(A[16]), .B(n30), .Z(n394) );
  GTECH_OAI21 U391 ( .A(n398), .B(n31), .C(n399), .Z(n397) );
  GTECH_OAI21 U392 ( .A(n266), .B(n305), .C(n400), .Z(n399) );
  GTECH_NOT U393 ( .A(n30), .Z(n299) );
  GTECH_NAND2 U394 ( .A(n282), .B(n401), .Z(N115) );
  GTECH_NOT U395 ( .A(N41), .Z(n401) );
  GTECH_NAND2 U396 ( .A(n289), .B(n283), .Z(N41) );
  GTECH_NAND2 U397 ( .A(Ld), .B(n289), .Z(n283) );
  GTECH_NOT U398 ( .A(n402), .Z(N113) );
  GTECH_AOI222 U399 ( .A(n271), .B(n305), .C(n273), .D(n306), .E(n304), .F(
        n269), .Z(n402) );
  GTECH_XOR2 U400 ( .A(n403), .B(n396), .Z(n304) );
  GTECH_ADD_ABC U401 ( .A(n32), .B(n265), .C(n404), .COUT(n396) );
  GTECH_NOT U402 ( .A(n405), .Z(n306) );
  GTECH_XOR2 U403 ( .A(n403), .B(n406), .Z(n405) );
  GTECH_NOT U404 ( .A(n400), .Z(n406) );
  GTECH_OAI21 U405 ( .A(n32), .B(n407), .C(n408), .Z(n400) );
  GTECH_OAI21 U406 ( .A(n265), .B(n310), .C(n409), .Z(n408) );
  GTECH_XOR2 U407 ( .A(n398), .B(n31), .Z(n403) );
  GTECH_NOT U408 ( .A(n266), .Z(n398) );
  GTECH_NOT U409 ( .A(n31), .Z(n305) );
  GTECH_NOT U410 ( .A(n410), .Z(N112) );
  GTECH_AOI222 U411 ( .A(n271), .B(n310), .C(n273), .D(n311), .E(n309), .F(
        n269), .Z(n410) );
  GTECH_XOR2 U412 ( .A(n411), .B(n404), .Z(n309) );
  GTECH_ADD_ABC U413 ( .A(n33), .B(n264), .C(n412), .COUT(n404) );
  GTECH_NOT U414 ( .A(n413), .Z(n311) );
  GTECH_XOR2 U415 ( .A(n411), .B(n414), .Z(n413) );
  GTECH_NOT U416 ( .A(n409), .Z(n414) );
  GTECH_OAI21 U417 ( .A(n33), .B(n415), .C(n416), .Z(n409) );
  GTECH_OAI21 U418 ( .A(n264), .B(n314), .C(n417), .Z(n416) );
  GTECH_XOR2 U419 ( .A(n407), .B(n32), .Z(n411) );
  GTECH_NOT U420 ( .A(n265), .Z(n407) );
  GTECH_NOT U421 ( .A(n32), .Z(n310) );
  GTECH_NOT U422 ( .A(n418), .Z(N111) );
  GTECH_AOI222 U423 ( .A(n271), .B(n314), .C(n273), .D(n315), .E(n313), .F(
        n269), .Z(n418) );
  GTECH_XOR2 U424 ( .A(n419), .B(n412), .Z(n313) );
  GTECH_ADD_ABC U425 ( .A(n34), .B(n263), .C(n420), .COUT(n412) );
  GTECH_NOT U426 ( .A(n421), .Z(n315) );
  GTECH_XOR2 U427 ( .A(n419), .B(n422), .Z(n421) );
  GTECH_NOT U428 ( .A(n417), .Z(n422) );
  GTECH_OAI21 U429 ( .A(n34), .B(n423), .C(n424), .Z(n417) );
  GTECH_OAI21 U430 ( .A(n263), .B(n318), .C(n425), .Z(n424) );
  GTECH_XOR2 U431 ( .A(n415), .B(n33), .Z(n419) );
  GTECH_NOT U432 ( .A(n264), .Z(n415) );
  GTECH_NOT U433 ( .A(n33), .Z(n314) );
  GTECH_NOT U434 ( .A(n426), .Z(N110) );
  GTECH_AOI222 U435 ( .A(n271), .B(n318), .C(n273), .D(n319), .E(n317), .F(
        n269), .Z(n426) );
  GTECH_XOR2 U436 ( .A(n427), .B(n420), .Z(n317) );
  GTECH_ADD_ABC U437 ( .A(n35), .B(n262), .C(n428), .COUT(n420) );
  GTECH_NOT U438 ( .A(n429), .Z(n319) );
  GTECH_XOR2 U439 ( .A(n427), .B(n430), .Z(n429) );
  GTECH_NOT U440 ( .A(n425), .Z(n430) );
  GTECH_OAI21 U441 ( .A(n35), .B(n431), .C(n432), .Z(n425) );
  GTECH_OAI21 U442 ( .A(n262), .B(n322), .C(n433), .Z(n432) );
  GTECH_XOR2 U443 ( .A(n423), .B(n34), .Z(n427) );
  GTECH_NOT U444 ( .A(n263), .Z(n423) );
  GTECH_NOT U445 ( .A(n34), .Z(n318) );
  GTECH_NOT U446 ( .A(n434), .Z(N109) );
  GTECH_AOI222 U447 ( .A(n271), .B(n322), .C(n273), .D(n323), .E(n321), .F(
        n269), .Z(n434) );
  GTECH_XOR2 U448 ( .A(n435), .B(n428), .Z(n321) );
  GTECH_ADD_ABC U449 ( .A(n36), .B(n261), .C(n436), .COUT(n428) );
  GTECH_NOT U450 ( .A(n437), .Z(n323) );
  GTECH_XOR2 U451 ( .A(n435), .B(n438), .Z(n437) );
  GTECH_NOT U452 ( .A(n433), .Z(n438) );
  GTECH_OAI21 U453 ( .A(n36), .B(n439), .C(n440), .Z(n433) );
  GTECH_OAI21 U454 ( .A(n261), .B(n326), .C(n441), .Z(n440) );
  GTECH_XOR2 U455 ( .A(n431), .B(n35), .Z(n435) );
  GTECH_NOT U456 ( .A(n262), .Z(n431) );
  GTECH_NOT U457 ( .A(n35), .Z(n322) );
  GTECH_NOT U458 ( .A(n442), .Z(N108) );
  GTECH_AOI222 U459 ( .A(n271), .B(n326), .C(n273), .D(n327), .E(n325), .F(
        n269), .Z(n442) );
  GTECH_XOR2 U460 ( .A(n443), .B(n436), .Z(n325) );
  GTECH_ADD_ABC U461 ( .A(n37), .B(n260), .C(n444), .COUT(n436) );
  GTECH_NOT U462 ( .A(n445), .Z(n327) );
  GTECH_XOR2 U463 ( .A(n443), .B(n446), .Z(n445) );
  GTECH_NOT U464 ( .A(n441), .Z(n446) );
  GTECH_OAI21 U465 ( .A(n37), .B(n447), .C(n448), .Z(n441) );
  GTECH_OAI21 U466 ( .A(n260), .B(n330), .C(n449), .Z(n448) );
  GTECH_XOR2 U467 ( .A(n439), .B(n36), .Z(n443) );
  GTECH_NOT U468 ( .A(n261), .Z(n439) );
  GTECH_NOT U469 ( .A(n36), .Z(n326) );
  GTECH_NOT U470 ( .A(n450), .Z(N107) );
  GTECH_AOI222 U471 ( .A(n271), .B(n330), .C(n273), .D(n331), .E(n329), .F(
        n269), .Z(n450) );
  GTECH_XOR2 U472 ( .A(n451), .B(n444), .Z(n329) );
  GTECH_ADD_ABC U473 ( .A(n38), .B(n259), .C(n452), .COUT(n444) );
  GTECH_NOT U474 ( .A(n453), .Z(n331) );
  GTECH_XOR2 U475 ( .A(n451), .B(n454), .Z(n453) );
  GTECH_NOT U476 ( .A(n449), .Z(n454) );
  GTECH_OAI21 U477 ( .A(n38), .B(n455), .C(n456), .Z(n449) );
  GTECH_OAI21 U478 ( .A(n259), .B(n334), .C(n457), .Z(n456) );
  GTECH_XOR2 U479 ( .A(n447), .B(n37), .Z(n451) );
  GTECH_NOT U480 ( .A(n260), .Z(n447) );
  GTECH_NOT U481 ( .A(n37), .Z(n330) );
  GTECH_NOT U482 ( .A(n458), .Z(N106) );
  GTECH_AOI222 U483 ( .A(n271), .B(n334), .C(n273), .D(n335), .E(n333), .F(
        n269), .Z(n458) );
  GTECH_XOR2 U484 ( .A(n459), .B(n452), .Z(n333) );
  GTECH_ADD_ABC U485 ( .A(n39), .B(n258), .C(n460), .COUT(n452) );
  GTECH_NOT U486 ( .A(n461), .Z(n335) );
  GTECH_XOR2 U487 ( .A(n459), .B(n462), .Z(n461) );
  GTECH_NOT U488 ( .A(n457), .Z(n462) );
  GTECH_OAI21 U489 ( .A(n39), .B(n463), .C(n464), .Z(n457) );
  GTECH_OAI21 U490 ( .A(n258), .B(n338), .C(n465), .Z(n464) );
  GTECH_XOR2 U491 ( .A(n455), .B(n38), .Z(n459) );
  GTECH_NOT U492 ( .A(n259), .Z(n455) );
  GTECH_NOT U493 ( .A(n38), .Z(n334) );
  GTECH_NOT U494 ( .A(n466), .Z(N105) );
  GTECH_AOI222 U495 ( .A(n271), .B(n338), .C(n273), .D(n339), .E(n337), .F(
        n269), .Z(n466) );
  GTECH_XOR2 U496 ( .A(n467), .B(n460), .Z(n337) );
  GTECH_ADD_ABC U497 ( .A(n40), .B(n257), .C(n468), .COUT(n460) );
  GTECH_NOT U498 ( .A(n469), .Z(n339) );
  GTECH_XOR2 U499 ( .A(n467), .B(n470), .Z(n469) );
  GTECH_NOT U500 ( .A(n465), .Z(n470) );
  GTECH_OAI21 U501 ( .A(n40), .B(n471), .C(n472), .Z(n465) );
  GTECH_OAI21 U502 ( .A(n257), .B(n342), .C(n473), .Z(n472) );
  GTECH_XOR2 U503 ( .A(n463), .B(n39), .Z(n467) );
  GTECH_NOT U504 ( .A(n258), .Z(n463) );
  GTECH_NOT U505 ( .A(n39), .Z(n338) );
  GTECH_NOT U506 ( .A(n474), .Z(N104) );
  GTECH_AOI222 U507 ( .A(n271), .B(n342), .C(n273), .D(n343), .E(n341), .F(
        n269), .Z(n474) );
  GTECH_XOR2 U508 ( .A(n475), .B(n468), .Z(n341) );
  GTECH_ADD_ABC U509 ( .A(n41), .B(n256), .C(n476), .COUT(n468) );
  GTECH_NOT U510 ( .A(n477), .Z(n343) );
  GTECH_XOR2 U511 ( .A(n475), .B(n478), .Z(n477) );
  GTECH_NOT U512 ( .A(n473), .Z(n478) );
  GTECH_OAI21 U513 ( .A(n41), .B(n479), .C(n480), .Z(n473) );
  GTECH_OAI21 U514 ( .A(n256), .B(n346), .C(n481), .Z(n480) );
  GTECH_XOR2 U515 ( .A(n471), .B(n40), .Z(n475) );
  GTECH_NOT U516 ( .A(n257), .Z(n471) );
  GTECH_NOT U517 ( .A(n40), .Z(n342) );
  GTECH_NOT U518 ( .A(n482), .Z(N103) );
  GTECH_AOI222 U519 ( .A(n271), .B(n346), .C(n273), .D(n347), .E(n345), .F(
        n269), .Z(n482) );
  GTECH_XOR2 U520 ( .A(n483), .B(n476), .Z(n345) );
  GTECH_ADD_ABC U521 ( .A(n42), .B(n255), .C(n484), .COUT(n476) );
  GTECH_NOT U522 ( .A(n485), .Z(n347) );
  GTECH_XOR2 U523 ( .A(n483), .B(n486), .Z(n485) );
  GTECH_NOT U524 ( .A(n481), .Z(n486) );
  GTECH_OAI21 U525 ( .A(n42), .B(n487), .C(n488), .Z(n481) );
  GTECH_OAI21 U526 ( .A(n255), .B(n351), .C(n489), .Z(n488) );
  GTECH_XOR2 U527 ( .A(n479), .B(n41), .Z(n483) );
  GTECH_NOT U528 ( .A(n256), .Z(n479) );
  GTECH_NOT U529 ( .A(n41), .Z(n346) );
  GTECH_NOT U530 ( .A(n490), .Z(N102) );
  GTECH_AOI222 U531 ( .A(n271), .B(n351), .C(n273), .D(n352), .E(n350), .F(
        n269), .Z(n490) );
  GTECH_XOR2 U532 ( .A(n491), .B(n484), .Z(n350) );
  GTECH_ADD_ABC U533 ( .A(n43), .B(n254), .C(n492), .COUT(n484) );
  GTECH_NOT U534 ( .A(n493), .Z(n352) );
  GTECH_XOR2 U535 ( .A(n491), .B(n494), .Z(n493) );
  GTECH_NOT U536 ( .A(n489), .Z(n494) );
  GTECH_OAI21 U537 ( .A(n43), .B(n495), .C(n496), .Z(n489) );
  GTECH_OAI21 U538 ( .A(n254), .B(n355), .C(n497), .Z(n496) );
  GTECH_XOR2 U539 ( .A(n487), .B(n42), .Z(n491) );
  GTECH_NOT U540 ( .A(n255), .Z(n487) );
  GTECH_NOT U541 ( .A(n42), .Z(n351) );
  GTECH_NOT U542 ( .A(n498), .Z(N101) );
  GTECH_AOI222 U543 ( .A(n271), .B(n355), .C(n273), .D(n356), .E(n354), .F(
        n269), .Z(n498) );
  GTECH_XOR2 U544 ( .A(n499), .B(n492), .Z(n354) );
  GTECH_ADD_ABC U545 ( .A(n29), .B(n253), .C(n500), .COUT(n492) );
  GTECH_NOT U546 ( .A(n501), .Z(n356) );
  GTECH_XOR2 U547 ( .A(n499), .B(n502), .Z(n501) );
  GTECH_NOT U548 ( .A(n497), .Z(n502) );
  GTECH_OAI21 U549 ( .A(n29), .B(n503), .C(n504), .Z(n497) );
  GTECH_OAI21 U550 ( .A(n253), .B(n359), .C(n505), .Z(n504) );
  GTECH_XOR2 U551 ( .A(n495), .B(n43), .Z(n499) );
  GTECH_NOT U552 ( .A(n254), .Z(n495) );
  GTECH_NOT U553 ( .A(n43), .Z(n355) );
  GTECH_NOT U554 ( .A(n506), .Z(N100) );
  GTECH_AOI222 U555 ( .A(n358), .B(n269), .C(n271), .D(n359), .E(n273), .F(
        n360), .Z(n506) );
  GTECH_NOT U556 ( .A(n507), .Z(n360) );
  GTECH_XOR2 U557 ( .A(n508), .B(n509), .Z(n507) );
  GTECH_NOT U558 ( .A(n505), .Z(n509) );
  GTECH_OAI21 U559 ( .A(n11), .B(n510), .C(n511), .Z(n505) );
  GTECH_OAI21 U560 ( .A(n252), .B(n272), .C(n365), .Z(n511) );
  GTECH_NAND2 U561 ( .A(n12), .B(n371), .Z(n365) );
  GTECH_NOT U562 ( .A(n11), .Z(n272) );
  GTECH_NOT U563 ( .A(n252), .Z(n510) );
  GTECH_NOT U564 ( .A(n281), .Z(n273) );
  GTECH_NAND2 U565 ( .A(N82), .B(n10), .Z(n281) );
  GTECH_NOT U566 ( .A(n512), .Z(N82) );
  GTECH_NOT U567 ( .A(n29), .Z(n359) );
  GTECH_NOT U568 ( .A(n513), .Z(n271) );
  GTECH_MUX2 U569 ( .A(n512), .B(n514), .S(n10), .Z(n513) );
  GTECH_NAND2 U570 ( .A(n28), .B(n287), .Z(n514) );
  GTECH_NAND2 U571 ( .A(n287), .B(n375), .Z(n512) );
  GTECH_NOT U572 ( .A(n28), .Z(n375) );
  GTECH_NOT U573 ( .A(n280), .Z(n269) );
  GTECH_NAND3 U574 ( .A(n287), .B(n373), .C(n28), .Z(n280) );
  GTECH_NOT U575 ( .A(n10), .Z(n373) );
  GTECH_NOT U576 ( .A(n282), .Z(n287) );
  GTECH_OAI21 U577 ( .A(n285), .B(n286), .C(n515), .Z(n282) );
  GTECH_AND2 U578 ( .A(n288), .B(n289), .Z(n515) );
  GTECH_NOT U579 ( .A(Rst), .Z(n289) );
  GTECH_NOT U580 ( .A(Ld), .Z(n288) );
  GTECH_NOT U581 ( .A(n9), .Z(n286) );
  GTECH_NAND2 U582 ( .A(n8), .B(n291), .Z(n285) );
  GTECH_NOT U583 ( .A(n294), .Z(n291) );
  GTECH_NAND2 U584 ( .A(n7), .B(n293), .Z(n294) );
  GTECH_NOT U585 ( .A(n516), .Z(n293) );
  GTECH_NAND2 U586 ( .A(n6), .B(n250), .Z(n516) );
  GTECH_XOR2 U587 ( .A(n508), .B(n500), .Z(n358) );
  GTECH_ADD_ABC U588 ( .A(n252), .B(n11), .C(n369), .COUT(n500) );
  GTECH_NAND2 U589 ( .A(n276), .B(n371), .Z(n369) );
  GTECH_NOT U590 ( .A(n251), .Z(n371) );
  GTECH_NOT U591 ( .A(n12), .Z(n276) );
  GTECH_XOR2 U592 ( .A(n503), .B(n29), .Z(n508) );
  GTECH_NOT U593 ( .A(n253), .Z(n503) );
endmodule

