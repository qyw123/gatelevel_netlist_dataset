
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130;

  GTECH_XOR2 U84 ( .A(n65), .B(n66), .Z(sum[9]) );
  GTECH_XNOR2 U85 ( .A(n67), .B(n68), .Z(sum[8]) );
  GTECH_XOR2 U86 ( .A(n69), .B(n70), .Z(sum[7]) );
  GTECH_OA21 U87 ( .A(n71), .B(n72), .C(n73), .Z(n70) );
  GTECH_XOR2 U88 ( .A(n72), .B(n71), .Z(sum[6]) );
  GTECH_OA21 U89 ( .A(n74), .B(n75), .C(n76), .Z(n71) );
  GTECH_XOR2 U90 ( .A(n75), .B(n74), .Z(sum[5]) );
  GTECH_OA21 U91 ( .A(n77), .B(n78), .C(n79), .Z(n74) );
  GTECH_XOR2 U92 ( .A(n78), .B(n77), .Z(sum[4]) );
  GTECH_XOR2 U93 ( .A(n80), .B(n81), .Z(sum[3]) );
  GTECH_OA21 U94 ( .A(n82), .B(n83), .C(n84), .Z(n81) );
  GTECH_XOR2 U95 ( .A(n82), .B(n83), .Z(sum[2]) );
  GTECH_AOI22 U96 ( .A(b[1]), .B(a[1]), .C(n85), .D(n86), .Z(n82) );
  GTECH_XOR2 U97 ( .A(n86), .B(n85), .Z(sum[1]) );
  GTECH_OAI2N2 U98 ( .A(n87), .B(n88), .C(a[0]), .D(b[0]), .Z(n85) );
  GTECH_XNOR2 U99 ( .A(n89), .B(n90), .Z(sum[15]) );
  GTECH_OAI21 U100 ( .A(n91), .B(n92), .C(n93), .Z(n89) );
  GTECH_XOR2 U101 ( .A(n92), .B(n91), .Z(sum[14]) );
  GTECH_OA21 U102 ( .A(n94), .B(n95), .C(n96), .Z(n91) );
  GTECH_XOR2 U103 ( .A(n95), .B(n94), .Z(sum[13]) );
  GTECH_OA21 U104 ( .A(n97), .B(n98), .C(n99), .Z(n94) );
  GTECH_NOT U105 ( .A(cout), .Z(n97) );
  GTECH_XNOR2 U106 ( .A(n98), .B(cout), .Z(sum[12]) );
  GTECH_XNOR2 U107 ( .A(n100), .B(n101), .Z(sum[11]) );
  GTECH_OAI21 U108 ( .A(n102), .B(n103), .C(n104), .Z(n100) );
  GTECH_XOR2 U109 ( .A(n103), .B(n102), .Z(sum[10]) );
  GTECH_OA21 U110 ( .A(n66), .B(n65), .C(n105), .Z(n102) );
  GTECH_OA21 U111 ( .A(n106), .B(n67), .C(n107), .Z(n66) );
  GTECH_NOT U112 ( .A(n68), .Z(n106) );
  GTECH_XNOR2 U113 ( .A(cin), .B(n87), .Z(sum[0]) );
  GTECH_AO21 U114 ( .A(n68), .B(n108), .C(n109), .Z(cout) );
  GTECH_OAI21 U115 ( .A(n77), .B(n110), .C(n111), .Z(n68) );
  GTECH_OA21 U116 ( .A(n112), .B(n88), .C(n113), .Z(n77) );
  GTECH_NOT U117 ( .A(cin), .Z(n88) );
  GTECH_NOR3 U118 ( .A(n110), .B(n112), .C(n114), .Z(Pm) );
  GTECH_OR5 U119 ( .A(n80), .B(n115), .C(n87), .D(n116), .E(n83), .Z(n112) );
  GTECH_XNOR2 U120 ( .A(a[0]), .B(b[0]), .Z(n87) );
  GTECH_AO21 U121 ( .A(n117), .B(n108), .C(n109), .Z(Gm) );
  GTECH_OAI21 U122 ( .A(n118), .B(n90), .C(n119), .Z(n109) );
  GTECH_OA21 U123 ( .A(n120), .B(n92), .C(n93), .Z(n118) );
  GTECH_OA21 U124 ( .A(n99), .B(n95), .C(n96), .Z(n120) );
  GTECH_NOT U125 ( .A(n114), .Z(n108) );
  GTECH_OR4 U126 ( .A(n98), .B(n90), .C(n92), .D(n95), .Z(n114) );
  GTECH_OAI21 U127 ( .A(b[13]), .B(a[13]), .C(n96), .Z(n95) );
  GTECH_NAND2 U128 ( .A(b[13]), .B(a[13]), .Z(n96) );
  GTECH_OAI21 U129 ( .A(b[14]), .B(a[14]), .C(n93), .Z(n92) );
  GTECH_NAND2 U130 ( .A(b[14]), .B(a[14]), .Z(n93) );
  GTECH_OAI21 U131 ( .A(b[15]), .B(a[15]), .C(n119), .Z(n90) );
  GTECH_NAND2 U132 ( .A(a[15]), .B(b[15]), .Z(n119) );
  GTECH_OAI21 U133 ( .A(b[12]), .B(a[12]), .C(n99), .Z(n98) );
  GTECH_NAND2 U134 ( .A(a[12]), .B(b[12]), .Z(n99) );
  GTECH_OAI21 U135 ( .A(n113), .B(n110), .C(n111), .Z(n117) );
  GTECH_OA21 U136 ( .A(n121), .B(n101), .C(n122), .Z(n111) );
  GTECH_OA21 U137 ( .A(n123), .B(n103), .C(n104), .Z(n121) );
  GTECH_OA21 U138 ( .A(n107), .B(n65), .C(n105), .Z(n123) );
  GTECH_OR4 U139 ( .A(n67), .B(n101), .C(n103), .D(n65), .Z(n110) );
  GTECH_OAI21 U140 ( .A(b[9]), .B(a[9]), .C(n105), .Z(n65) );
  GTECH_NAND2 U141 ( .A(a[9]), .B(b[9]), .Z(n105) );
  GTECH_OAI21 U142 ( .A(b[10]), .B(a[10]), .C(n104), .Z(n103) );
  GTECH_NAND2 U143 ( .A(b[10]), .B(a[10]), .Z(n104) );
  GTECH_OAI21 U144 ( .A(b[11]), .B(a[11]), .C(n122), .Z(n101) );
  GTECH_NAND2 U145 ( .A(a[11]), .B(b[11]), .Z(n122) );
  GTECH_OAI21 U146 ( .A(b[8]), .B(a[8]), .C(n107), .Z(n67) );
  GTECH_NAND2 U147 ( .A(a[8]), .B(b[8]), .Z(n107) );
  GTECH_AOI21 U148 ( .A(b[7]), .B(a[7]), .C(n124), .Z(n113) );
  GTECH_OAI22 U149 ( .A(n125), .B(n116), .C(n126), .D(n69), .Z(n124) );
  GTECH_OA21 U150 ( .A(n127), .B(n72), .C(n73), .Z(n126) );
  GTECH_OA21 U151 ( .A(n75), .B(n79), .C(n76), .Z(n127) );
  GTECH_OR4 U152 ( .A(n75), .B(n72), .C(n78), .D(n69), .Z(n116) );
  GTECH_XNOR2 U153 ( .A(a[7]), .B(b[7]), .Z(n69) );
  GTECH_OAI21 U154 ( .A(b[4]), .B(a[4]), .C(n79), .Z(n78) );
  GTECH_NAND2 U155 ( .A(b[4]), .B(a[4]), .Z(n79) );
  GTECH_OAI21 U156 ( .A(b[6]), .B(a[6]), .C(n73), .Z(n72) );
  GTECH_NAND2 U157 ( .A(b[6]), .B(a[6]), .Z(n73) );
  GTECH_OAI21 U158 ( .A(b[5]), .B(a[5]), .C(n76), .Z(n75) );
  GTECH_NAND2 U159 ( .A(b[5]), .B(a[5]), .Z(n76) );
  GTECH_AOI2N2 U160 ( .A(b[3]), .B(a[3]), .C(n128), .D(n80), .Z(n125) );
  GTECH_XNOR2 U161 ( .A(a[3]), .B(b[3]), .Z(n80) );
  GTECH_OA21 U162 ( .A(n129), .B(n83), .C(n84), .Z(n128) );
  GTECH_OAI21 U163 ( .A(a[2]), .B(b[2]), .C(n84), .Z(n83) );
  GTECH_NAND2 U164 ( .A(b[2]), .B(a[2]), .Z(n84) );
  GTECH_AOI21 U165 ( .A(b[1]), .B(a[1]), .C(n130), .Z(n129) );
  GTECH_AND3 U166 ( .A(a[0]), .B(n86), .C(b[0]), .Z(n130) );
  GTECH_NOT U167 ( .A(n115), .Z(n86) );
  GTECH_XNOR2 U168 ( .A(a[1]), .B(b[1]), .Z(n115) );
endmodule

