
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_OR_NOT U83 ( .A(n97), .B(n93), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n98), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n98) );
  GTECH_OAI21 U86 ( .A(n99), .B(n100), .C(n101), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  GTECH_NOT U88 ( .A(n103), .Z(n99) );
  GTECH_OR_NOT U89 ( .A(n105), .B(I_b[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n106), .Z(n84) );
  GTECH_OR_NOT U91 ( .A(n107), .B(n108), .Z(n106) );
  GTECH_XOR2 U92 ( .A(n109), .B(n108), .Z(N153) );
  GTECH_NOT U93 ( .A(n110), .Z(n108) );
  GTECH_XOR3 U94 ( .A(n97), .B(n93), .C(n95), .Z(n110) );
  GTECH_XOR3 U95 ( .A(n102), .B(n104), .C(n103), .Z(n95) );
  GTECH_OAI21 U96 ( .A(n111), .B(n112), .C(n113), .Z(n103) );
  GTECH_OAI21 U97 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_NOT U98 ( .A(n115), .Z(n111) );
  GTECH_NOT U99 ( .A(n117), .Z(n104) );
  GTECH_OR_NOT U100 ( .A(n118), .B(I_b[7]), .Z(n117) );
  GTECH_NOT U101 ( .A(n100), .Z(n102) );
  GTECH_OR_NOT U102 ( .A(n119), .B(I_a[7]), .Z(n100) );
  GTECH_NOT U103 ( .A(I_b[6]), .Z(n119) );
  GTECH_ADD_ABC U104 ( .A(n120), .B(n121), .C(n122), .COUT(n93) );
  GTECH_NOT U105 ( .A(n123), .Z(n122) );
  GTECH_XOR2 U106 ( .A(n124), .B(n125), .Z(n121) );
  GTECH_AND_NOT U107 ( .A(I_a[7]), .B(n126), .Z(n125) );
  GTECH_NOT U108 ( .A(n94), .Z(n97) );
  GTECH_OR_NOT U109 ( .A(n124), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U110 ( .A(n107), .Z(n109) );
  GTECH_OR_NOT U111 ( .A(n127), .B(n128), .Z(n107) );
  GTECH_XOR2 U112 ( .A(n127), .B(n129), .Z(N152) );
  GTECH_NOT U113 ( .A(n128), .Z(n129) );
  GTECH_XOR4 U114 ( .A(n130), .B(n124), .C(n120), .D(n123), .Z(n128) );
  GTECH_XOR3 U115 ( .A(n114), .B(n116), .C(n115), .Z(n123) );
  GTECH_OAI21 U116 ( .A(n131), .B(n132), .C(n133), .Z(n115) );
  GTECH_OAI21 U117 ( .A(n134), .B(n135), .C(n136), .Z(n133) );
  GTECH_NOT U118 ( .A(n135), .Z(n131) );
  GTECH_NOT U119 ( .A(n137), .Z(n116) );
  GTECH_OR_NOT U120 ( .A(n138), .B(I_b[7]), .Z(n137) );
  GTECH_NOT U121 ( .A(n112), .Z(n114) );
  GTECH_OR_NOT U122 ( .A(n118), .B(I_b[6]), .Z(n112) );
  GTECH_NOT U123 ( .A(I_a[6]), .Z(n118) );
  GTECH_ADD_ABC U124 ( .A(n139), .B(n140), .C(n141), .COUT(n120) );
  GTECH_NOT U125 ( .A(n142), .Z(n141) );
  GTECH_XOR3 U126 ( .A(n143), .B(n144), .C(n145), .Z(n140) );
  GTECH_OA21 U127 ( .A(n145), .B(n146), .C(n147), .Z(n124) );
  GTECH_OAI21 U128 ( .A(n143), .B(n148), .C(n144), .Z(n147) );
  GTECH_NOT U129 ( .A(n146), .Z(n143) );
  GTECH_NOT U130 ( .A(n148), .Z(n145) );
  GTECH_AND_NOT U131 ( .A(I_a[7]), .B(n126), .Z(n130) );
  GTECH_ADD_ABC U132 ( .A(n149), .B(n150), .C(n151), .COUT(n127) );
  GTECH_NOT U133 ( .A(n152), .Z(n151) );
  GTECH_OA22 U134 ( .A(n153), .B(n105), .C(n154), .D(n155), .Z(n150) );
  GTECH_OA21 U135 ( .A(n156), .B(n157), .C(n158), .Z(n149) );
  GTECH_XOR3 U136 ( .A(n159), .B(n152), .C(n160), .Z(N151) );
  GTECH_OA21 U137 ( .A(n156), .B(n157), .C(n158), .Z(n160) );
  GTECH_OAI21 U138 ( .A(n161), .B(n162), .C(n163), .Z(n158) );
  GTECH_XOR2 U139 ( .A(n164), .B(n139), .Z(n152) );
  GTECH_ADD_ABC U140 ( .A(n165), .B(n166), .C(n167), .COUT(n139) );
  GTECH_NOT U141 ( .A(n168), .Z(n167) );
  GTECH_XOR3 U142 ( .A(n169), .B(n170), .C(n171), .Z(n166) );
  GTECH_XOR4 U143 ( .A(n144), .B(n148), .C(n146), .D(n142), .Z(n164) );
  GTECH_XOR3 U144 ( .A(n134), .B(n136), .C(n135), .Z(n142) );
  GTECH_OAI21 U145 ( .A(n172), .B(n173), .C(n174), .Z(n135) );
  GTECH_OAI21 U146 ( .A(n175), .B(n176), .C(n177), .Z(n174) );
  GTECH_NOT U147 ( .A(n176), .Z(n172) );
  GTECH_NOT U148 ( .A(n178), .Z(n136) );
  GTECH_OR_NOT U149 ( .A(n179), .B(I_b[7]), .Z(n178) );
  GTECH_NOT U150 ( .A(n132), .Z(n134) );
  GTECH_OR_NOT U151 ( .A(n138), .B(I_b[6]), .Z(n132) );
  GTECH_NOT U152 ( .A(I_a[5]), .Z(n138) );
  GTECH_OR_NOT U153 ( .A(n180), .B(I_a[7]), .Z(n146) );
  GTECH_OAI21 U154 ( .A(n171), .B(n181), .C(n182), .Z(n148) );
  GTECH_OAI21 U155 ( .A(n169), .B(n183), .C(n170), .Z(n182) );
  GTECH_NOT U156 ( .A(n181), .Z(n169) );
  GTECH_NOT U157 ( .A(n183), .Z(n171) );
  GTECH_NOT U158 ( .A(n184), .Z(n144) );
  GTECH_OR_NOT U159 ( .A(n126), .B(I_a[6]), .Z(n184) );
  GTECH_OA22 U160 ( .A(n153), .B(n105), .C(n154), .D(n155), .Z(n159) );
  GTECH_NOT U161 ( .A(n185), .Z(n155) );
  GTECH_NOT U162 ( .A(I_a[7]), .Z(n105) );
  GTECH_XOR3 U163 ( .A(n156), .B(n161), .C(n186), .Z(N150) );
  GTECH_NOT U164 ( .A(n163), .Z(n186) );
  GTECH_XOR2 U165 ( .A(n187), .B(n165), .Z(n163) );
  GTECH_ADD_ABC U166 ( .A(n188), .B(n189), .C(n190), .COUT(n165) );
  GTECH_NOT U167 ( .A(n191), .Z(n190) );
  GTECH_XOR3 U168 ( .A(n192), .B(n193), .C(n194), .Z(n189) );
  GTECH_XOR4 U169 ( .A(n170), .B(n183), .C(n181), .D(n168), .Z(n187) );
  GTECH_XOR3 U170 ( .A(n175), .B(n177), .C(n176), .Z(n168) );
  GTECH_OAI21 U171 ( .A(n195), .B(n196), .C(n197), .Z(n176) );
  GTECH_OAI21 U172 ( .A(n198), .B(n199), .C(n200), .Z(n197) );
  GTECH_NOT U173 ( .A(n199), .Z(n195) );
  GTECH_NOT U174 ( .A(n201), .Z(n177) );
  GTECH_OR_NOT U175 ( .A(n202), .B(I_b[7]), .Z(n201) );
  GTECH_NOT U176 ( .A(n173), .Z(n175) );
  GTECH_OR_NOT U177 ( .A(n179), .B(I_b[6]), .Z(n173) );
  GTECH_OR_NOT U178 ( .A(n180), .B(I_a[6]), .Z(n181) );
  GTECH_OAI21 U179 ( .A(n194), .B(n203), .C(n204), .Z(n183) );
  GTECH_OAI21 U180 ( .A(n192), .B(n205), .C(n193), .Z(n204) );
  GTECH_NOT U181 ( .A(n203), .Z(n192) );
  GTECH_NOT U182 ( .A(n205), .Z(n194) );
  GTECH_NOT U183 ( .A(n206), .Z(n170) );
  GTECH_OR_NOT U184 ( .A(n126), .B(I_a[5]), .Z(n206) );
  GTECH_NOT U185 ( .A(I_b[5]), .Z(n126) );
  GTECH_NOT U186 ( .A(n157), .Z(n161) );
  GTECH_XOR2 U187 ( .A(n185), .B(n154), .Z(n157) );
  GTECH_AOI2N2 U188 ( .A(n207), .B(n208), .C(n209), .D(n210), .Z(n154) );
  GTECH_OR_NOT U189 ( .A(n211), .B(n209), .Z(n208) );
  GTECH_XOR2 U190 ( .A(n212), .B(n153), .Z(n185) );
  GTECH_OA21 U191 ( .A(n213), .B(n214), .C(n215), .Z(n153) );
  GTECH_OR_NOT U192 ( .A(n216), .B(n217), .Z(n215) );
  GTECH_AND_NOT U193 ( .A(n216), .B(n217), .Z(n213) );
  GTECH_OR_NOT U194 ( .A(n218), .B(I_a[7]), .Z(n212) );
  GTECH_NOT U195 ( .A(n162), .Z(n156) );
  GTECH_OAI2N2 U196 ( .A(n219), .B(n220), .C(n221), .D(n222), .Z(n162) );
  GTECH_OR_NOT U197 ( .A(n223), .B(n219), .Z(n222) );
  GTECH_XOR3 U198 ( .A(n219), .B(n223), .C(n224), .Z(N149) );
  GTECH_NOT U199 ( .A(n221), .Z(n224) );
  GTECH_XOR2 U200 ( .A(n225), .B(n188), .Z(n221) );
  GTECH_ADD_ABC U201 ( .A(n226), .B(n227), .C(n228), .COUT(n188) );
  GTECH_XOR3 U202 ( .A(n229), .B(n230), .C(n231), .Z(n227) );
  GTECH_OA21 U203 ( .A(n232), .B(n233), .C(n234), .Z(n226) );
  GTECH_XOR4 U204 ( .A(n193), .B(n205), .C(n203), .D(n191), .Z(n225) );
  GTECH_XOR3 U205 ( .A(n198), .B(n200), .C(n199), .Z(n191) );
  GTECH_OAI21 U206 ( .A(n235), .B(n236), .C(n237), .Z(n199) );
  GTECH_NOT U207 ( .A(n238), .Z(n200) );
  GTECH_OR_NOT U208 ( .A(n239), .B(I_b[7]), .Z(n238) );
  GTECH_NOT U209 ( .A(n196), .Z(n198) );
  GTECH_OR_NOT U210 ( .A(n202), .B(I_b[6]), .Z(n196) );
  GTECH_OR_NOT U211 ( .A(n180), .B(I_a[5]), .Z(n203) );
  GTECH_NOT U212 ( .A(I_b[4]), .Z(n180) );
  GTECH_OAI21 U213 ( .A(n231), .B(n240), .C(n241), .Z(n205) );
  GTECH_OAI21 U214 ( .A(n229), .B(n242), .C(n230), .Z(n241) );
  GTECH_NOT U215 ( .A(n240), .Z(n229) );
  GTECH_NOT U216 ( .A(n242), .Z(n231) );
  GTECH_NOT U217 ( .A(n243), .Z(n193) );
  GTECH_OR_NOT U218 ( .A(n179), .B(I_b[5]), .Z(n243) );
  GTECH_NOT U219 ( .A(n220), .Z(n223) );
  GTECH_XOR3 U220 ( .A(n211), .B(n209), .C(n207), .Z(n220) );
  GTECH_XOR3 U221 ( .A(n244), .B(n245), .C(n217), .Z(n207) );
  GTECH_OAI21 U222 ( .A(n246), .B(n247), .C(n248), .Z(n217) );
  GTECH_OAI21 U223 ( .A(n249), .B(n250), .C(n251), .Z(n248) );
  GTECH_NOT U224 ( .A(n250), .Z(n246) );
  GTECH_NOT U225 ( .A(n214), .Z(n245) );
  GTECH_OR_NOT U226 ( .A(n218), .B(I_a[6]), .Z(n214) );
  GTECH_NOT U227 ( .A(n216), .Z(n244) );
  GTECH_OR_NOT U228 ( .A(n252), .B(I_a[7]), .Z(n216) );
  GTECH_ADD_ABC U229 ( .A(n253), .B(n254), .C(n255), .COUT(n209) );
  GTECH_XOR2 U230 ( .A(n256), .B(n257), .Z(n254) );
  GTECH_AND_NOT U231 ( .A(I_a[7]), .B(n258), .Z(n257) );
  GTECH_NOT U232 ( .A(n210), .Z(n211) );
  GTECH_OR_NOT U233 ( .A(n256), .B(I_a[7]), .Z(n210) );
  GTECH_ADD_ABC U234 ( .A(n259), .B(n260), .C(n261), .COUT(n219) );
  GTECH_XOR3 U235 ( .A(n253), .B(n262), .C(n255), .Z(n260) );
  GTECH_NOT U236 ( .A(n263), .Z(n255) );
  GTECH_XOR2 U237 ( .A(n259), .B(n264), .Z(N148) );
  GTECH_XOR4 U238 ( .A(n262), .B(n263), .C(n261), .D(n253), .Z(n264) );
  GTECH_ADD_ABC U239 ( .A(n265), .B(n266), .C(n267), .COUT(n253) );
  GTECH_XOR3 U240 ( .A(n268), .B(n269), .C(n270), .Z(n266) );
  GTECH_XOR2 U241 ( .A(n271), .B(n272), .Z(n261) );
  GTECH_OA21 U242 ( .A(n232), .B(n233), .C(n234), .Z(n272) );
  GTECH_OAI21 U243 ( .A(n273), .B(n274), .C(n275), .Z(n234) );
  GTECH_NOT U244 ( .A(n232), .Z(n274) );
  GTECH_XOR4 U245 ( .A(n230), .B(n242), .C(n240), .D(n228), .Z(n271) );
  GTECH_XOR3 U246 ( .A(n276), .B(n277), .C(n237), .Z(n228) );
  GTECH_NAND3 U247 ( .A(I_b[6]), .B(I_a[1]), .C(n278), .Z(n237) );
  GTECH_NOT U248 ( .A(n236), .Z(n277) );
  GTECH_OR_NOT U249 ( .A(n279), .B(I_b[7]), .Z(n236) );
  GTECH_NOT U250 ( .A(n235), .Z(n276) );
  GTECH_OR_NOT U251 ( .A(n239), .B(I_b[6]), .Z(n235) );
  GTECH_OR_NOT U252 ( .A(n179), .B(I_b[4]), .Z(n240) );
  GTECH_OAI21 U253 ( .A(n280), .B(n281), .C(n282), .Z(n242) );
  GTECH_OAI21 U254 ( .A(n283), .B(n284), .C(n285), .Z(n282) );
  GTECH_NOT U255 ( .A(n284), .Z(n280) );
  GTECH_NOT U256 ( .A(n286), .Z(n230) );
  GTECH_OR_NOT U257 ( .A(n202), .B(I_b[5]), .Z(n286) );
  GTECH_XOR3 U258 ( .A(n249), .B(n251), .C(n250), .Z(n263) );
  GTECH_OAI21 U259 ( .A(n287), .B(n288), .C(n289), .Z(n250) );
  GTECH_OAI21 U260 ( .A(n290), .B(n291), .C(n292), .Z(n289) );
  GTECH_NOT U261 ( .A(n291), .Z(n287) );
  GTECH_NOT U262 ( .A(n293), .Z(n251) );
  GTECH_OR_NOT U263 ( .A(n218), .B(I_a[5]), .Z(n293) );
  GTECH_NOT U264 ( .A(I_b[3]), .Z(n218) );
  GTECH_NOT U265 ( .A(n247), .Z(n249) );
  GTECH_OR_NOT U266 ( .A(n252), .B(I_a[6]), .Z(n247) );
  GTECH_XOR2 U267 ( .A(n294), .B(n256), .Z(n262) );
  GTECH_OA21 U268 ( .A(n270), .B(n295), .C(n296), .Z(n256) );
  GTECH_OAI21 U269 ( .A(n268), .B(n297), .C(n269), .Z(n296) );
  GTECH_NOT U270 ( .A(n297), .Z(n270) );
  GTECH_AND_NOT U271 ( .A(I_a[7]), .B(n258), .Z(n294) );
  GTECH_ADD_ABC U272 ( .A(n298), .B(n299), .C(n300), .COUT(n259) );
  GTECH_NOT U273 ( .A(n301), .Z(n300) );
  GTECH_XOR3 U274 ( .A(n265), .B(n302), .C(n267), .Z(n299) );
  GTECH_NOT U275 ( .A(n303), .Z(n267) );
  GTECH_NOT U276 ( .A(n304), .Z(n302) );
  GTECH_XOR2 U277 ( .A(n305), .B(n298), .Z(N147) );
  GTECH_ADD_ABC U278 ( .A(n306), .B(n307), .C(n308), .COUT(n298) );
  GTECH_XOR3 U279 ( .A(n309), .B(n310), .C(n311), .Z(n307) );
  GTECH_OA21 U280 ( .A(n312), .B(n313), .C(n314), .Z(n306) );
  GTECH_XOR4 U281 ( .A(n303), .B(n265), .C(n304), .D(n301), .Z(n305) );
  GTECH_XOR3 U282 ( .A(n275), .B(n233), .C(n232), .Z(n301) );
  GTECH_XOR2 U283 ( .A(n315), .B(n278), .Z(n232) );
  GTECH_NOT U284 ( .A(n316), .Z(n278) );
  GTECH_OR_NOT U285 ( .A(n317), .B(I_b[7]), .Z(n316) );
  GTECH_OR_NOT U286 ( .A(n279), .B(I_b[6]), .Z(n315) );
  GTECH_NOT U287 ( .A(n273), .Z(n233) );
  GTECH_XOR3 U288 ( .A(n283), .B(n285), .C(n284), .Z(n273) );
  GTECH_OAI21 U289 ( .A(n318), .B(n319), .C(n320), .Z(n284) );
  GTECH_NOT U290 ( .A(n321), .Z(n285) );
  GTECH_OR_NOT U291 ( .A(n239), .B(I_b[5]), .Z(n321) );
  GTECH_NOT U292 ( .A(n281), .Z(n283) );
  GTECH_OR_NOT U293 ( .A(n202), .B(I_b[4]), .Z(n281) );
  GTECH_NOT U294 ( .A(n322), .Z(n275) );
  GTECH_NAND3 U295 ( .A(I_a[0]), .B(n323), .C(I_b[6]), .Z(n322) );
  GTECH_NOT U296 ( .A(n324), .Z(n323) );
  GTECH_XOR3 U297 ( .A(n268), .B(n269), .C(n297), .Z(n304) );
  GTECH_OAI21 U298 ( .A(n325), .B(n326), .C(n327), .Z(n297) );
  GTECH_OAI21 U299 ( .A(n328), .B(n329), .C(n330), .Z(n327) );
  GTECH_NOT U300 ( .A(n331), .Z(n269) );
  GTECH_OR_NOT U301 ( .A(n258), .B(I_a[6]), .Z(n331) );
  GTECH_NOT U302 ( .A(n295), .Z(n268) );
  GTECH_OR_NOT U303 ( .A(n332), .B(I_a[7]), .Z(n295) );
  GTECH_ADD_ABC U304 ( .A(n309), .B(n333), .C(n311), .COUT(n265) );
  GTECH_NOT U305 ( .A(n334), .Z(n311) );
  GTECH_XOR3 U306 ( .A(n328), .B(n330), .C(n325), .Z(n333) );
  GTECH_NOT U307 ( .A(n329), .Z(n325) );
  GTECH_XOR3 U308 ( .A(n290), .B(n292), .C(n291), .Z(n303) );
  GTECH_OAI21 U309 ( .A(n335), .B(n336), .C(n337), .Z(n291) );
  GTECH_OAI21 U310 ( .A(n338), .B(n339), .C(n340), .Z(n337) );
  GTECH_NOT U311 ( .A(n339), .Z(n335) );
  GTECH_NOT U312 ( .A(n341), .Z(n292) );
  GTECH_OR_NOT U313 ( .A(n179), .B(I_b[3]), .Z(n341) );
  GTECH_NOT U314 ( .A(n288), .Z(n290) );
  GTECH_OR_NOT U315 ( .A(n252), .B(I_a[5]), .Z(n288) );
  GTECH_NOT U316 ( .A(I_b[2]), .Z(n252) );
  GTECH_XOR2 U317 ( .A(n342), .B(n343), .Z(N146) );
  GTECH_XOR4 U318 ( .A(n310), .B(n334), .C(n308), .D(n309), .Z(n343) );
  GTECH_ADD_ABC U319 ( .A(n344), .B(n345), .C(n346), .COUT(n309) );
  GTECH_NOT U320 ( .A(n347), .Z(n346) );
  GTECH_XOR3 U321 ( .A(n348), .B(n349), .C(n350), .Z(n345) );
  GTECH_XOR2 U322 ( .A(n324), .B(n351), .Z(n308) );
  GTECH_AND_NOT U323 ( .A(I_b[6]), .B(n317), .Z(n351) );
  GTECH_XOR3 U324 ( .A(n352), .B(n353), .C(n320), .Z(n324) );
  GTECH_NAND3 U325 ( .A(I_b[4]), .B(I_a[1]), .C(n354), .Z(n320) );
  GTECH_NOT U326 ( .A(n319), .Z(n353) );
  GTECH_OR_NOT U327 ( .A(n279), .B(I_b[5]), .Z(n319) );
  GTECH_NOT U328 ( .A(n318), .Z(n352) );
  GTECH_OR_NOT U329 ( .A(n239), .B(I_b[4]), .Z(n318) );
  GTECH_XOR3 U330 ( .A(n338), .B(n340), .C(n339), .Z(n334) );
  GTECH_OAI21 U331 ( .A(n355), .B(n356), .C(n357), .Z(n339) );
  GTECH_OAI21 U332 ( .A(n358), .B(n359), .C(n360), .Z(n357) );
  GTECH_NOT U333 ( .A(n359), .Z(n355) );
  GTECH_NOT U334 ( .A(n361), .Z(n340) );
  GTECH_OR_NOT U335 ( .A(n202), .B(I_b[3]), .Z(n361) );
  GTECH_NOT U336 ( .A(n336), .Z(n338) );
  GTECH_OR_NOT U337 ( .A(n179), .B(I_b[2]), .Z(n336) );
  GTECH_NOT U338 ( .A(I_a[4]), .Z(n179) );
  GTECH_NOT U339 ( .A(n362), .Z(n310) );
  GTECH_XOR3 U340 ( .A(n328), .B(n330), .C(n329), .Z(n362) );
  GTECH_OAI21 U341 ( .A(n350), .B(n363), .C(n364), .Z(n329) );
  GTECH_OAI21 U342 ( .A(n348), .B(n365), .C(n349), .Z(n364) );
  GTECH_NOT U343 ( .A(n363), .Z(n348) );
  GTECH_NOT U344 ( .A(n365), .Z(n350) );
  GTECH_NOT U345 ( .A(n366), .Z(n330) );
  GTECH_OR_NOT U346 ( .A(n258), .B(I_a[5]), .Z(n366) );
  GTECH_NOT U347 ( .A(n326), .Z(n328) );
  GTECH_OR_NOT U348 ( .A(n332), .B(I_a[6]), .Z(n326) );
  GTECH_OA21 U349 ( .A(n312), .B(n313), .C(n314), .Z(n342) );
  GTECH_OAI21 U350 ( .A(n367), .B(n368), .C(n369), .Z(n314) );
  GTECH_NOT U351 ( .A(n312), .Z(n368) );
  GTECH_XOR3 U352 ( .A(n369), .B(n313), .C(n312), .Z(N145) );
  GTECH_XOR2 U353 ( .A(n370), .B(n354), .Z(n312) );
  GTECH_NOT U354 ( .A(n371), .Z(n354) );
  GTECH_OR_NOT U355 ( .A(n317), .B(I_b[5]), .Z(n371) );
  GTECH_OR_NOT U356 ( .A(n279), .B(I_b[4]), .Z(n370) );
  GTECH_NOT U357 ( .A(n367), .Z(n313) );
  GTECH_XOR2 U358 ( .A(n372), .B(n344), .Z(n367) );
  GTECH_ADD_ABC U359 ( .A(n373), .B(n374), .C(n375), .COUT(n344) );
  GTECH_XOR3 U360 ( .A(n376), .B(n377), .C(n378), .Z(n374) );
  GTECH_OA21 U361 ( .A(n379), .B(n380), .C(n381), .Z(n373) );
  GTECH_XOR4 U362 ( .A(n349), .B(n365), .C(n363), .D(n347), .Z(n372) );
  GTECH_XOR3 U363 ( .A(n358), .B(n360), .C(n359), .Z(n347) );
  GTECH_OAI21 U364 ( .A(n382), .B(n383), .C(n384), .Z(n359) );
  GTECH_NOT U365 ( .A(n385), .Z(n360) );
  GTECH_OR_NOT U366 ( .A(n239), .B(I_b[3]), .Z(n385) );
  GTECH_NOT U367 ( .A(n356), .Z(n358) );
  GTECH_OR_NOT U368 ( .A(n202), .B(I_b[2]), .Z(n356) );
  GTECH_OR_NOT U369 ( .A(n332), .B(I_a[5]), .Z(n363) );
  GTECH_OAI21 U370 ( .A(n378), .B(n386), .C(n387), .Z(n365) );
  GTECH_OAI21 U371 ( .A(n376), .B(n388), .C(n377), .Z(n387) );
  GTECH_NOT U372 ( .A(n388), .Z(n378) );
  GTECH_NOT U373 ( .A(n389), .Z(n349) );
  GTECH_OR_NOT U374 ( .A(n258), .B(I_a[4]), .Z(n389) );
  GTECH_NOT U375 ( .A(n390), .Z(n369) );
  GTECH_NAND3 U376 ( .A(I_a[0]), .B(n391), .C(I_b[4]), .Z(n390) );
  GTECH_XOR2 U377 ( .A(n392), .B(n391), .Z(N144) );
  GTECH_XOR2 U378 ( .A(n393), .B(n394), .Z(n391) );
  GTECH_XOR4 U379 ( .A(n377), .B(n388), .C(n375), .D(n376), .Z(n394) );
  GTECH_NOT U380 ( .A(n386), .Z(n376) );
  GTECH_OR_NOT U381 ( .A(n332), .B(I_a[4]), .Z(n386) );
  GTECH_XOR3 U382 ( .A(n395), .B(n396), .C(n384), .Z(n375) );
  GTECH_NAND3 U383 ( .A(I_b[2]), .B(I_a[1]), .C(n397), .Z(n384) );
  GTECH_NOT U384 ( .A(n383), .Z(n396) );
  GTECH_OR_NOT U385 ( .A(n279), .B(I_b[3]), .Z(n383) );
  GTECH_NOT U386 ( .A(n382), .Z(n395) );
  GTECH_OR_NOT U387 ( .A(n239), .B(I_b[2]), .Z(n382) );
  GTECH_OAI21 U388 ( .A(n398), .B(n399), .C(n400), .Z(n388) );
  GTECH_OAI21 U389 ( .A(n401), .B(n402), .C(n403), .Z(n400) );
  GTECH_NOT U390 ( .A(n402), .Z(n398) );
  GTECH_NOT U391 ( .A(n404), .Z(n377) );
  GTECH_OR_NOT U392 ( .A(n258), .B(I_a[3]), .Z(n404) );
  GTECH_OA21 U393 ( .A(n379), .B(n380), .C(n381), .Z(n393) );
  GTECH_OAI21 U394 ( .A(n405), .B(n406), .C(n407), .Z(n381) );
  GTECH_NOT U395 ( .A(n379), .Z(n406) );
  GTECH_AND_NOT U396 ( .A(I_b[4]), .B(n317), .Z(n392) );
  GTECH_XOR3 U397 ( .A(n407), .B(n380), .C(n379), .Z(N143) );
  GTECH_XOR2 U398 ( .A(n408), .B(n397), .Z(n379) );
  GTECH_NOT U399 ( .A(n409), .Z(n397) );
  GTECH_OR_NOT U400 ( .A(n317), .B(I_b[3]), .Z(n409) );
  GTECH_OR_NOT U401 ( .A(n279), .B(I_b[2]), .Z(n408) );
  GTECH_NOT U402 ( .A(I_a[1]), .Z(n279) );
  GTECH_NOT U403 ( .A(n405), .Z(n380) );
  GTECH_XOR3 U404 ( .A(n401), .B(n403), .C(n402), .Z(n405) );
  GTECH_OAI21 U405 ( .A(n410), .B(n411), .C(n412), .Z(n402) );
  GTECH_NOT U406 ( .A(n413), .Z(n403) );
  GTECH_OR_NOT U407 ( .A(n239), .B(I_b[1]), .Z(n413) );
  GTECH_NOT U408 ( .A(n399), .Z(n401) );
  GTECH_OR_NOT U409 ( .A(n202), .B(I_b[0]), .Z(n399) );
  GTECH_NOT U410 ( .A(I_a[3]), .Z(n202) );
  GTECH_NOT U411 ( .A(n414), .Z(n407) );
  GTECH_NAND3 U412 ( .A(I_a[0]), .B(n415), .C(I_b[2]), .Z(n414) );
  GTECH_XOR2 U413 ( .A(n416), .B(n415), .Z(N142) );
  GTECH_NOT U414 ( .A(n417), .Z(n415) );
  GTECH_XOR3 U415 ( .A(n418), .B(n419), .C(n412), .Z(n417) );
  GTECH_NAND3 U416 ( .A(n420), .B(I_b[0]), .C(I_a[1]), .Z(n412) );
  GTECH_NOT U417 ( .A(n410), .Z(n419) );
  GTECH_OR_NOT U418 ( .A(n258), .B(I_a[1]), .Z(n410) );
  GTECH_NOT U419 ( .A(n411), .Z(n418) );
  GTECH_OR_NOT U420 ( .A(n239), .B(I_b[0]), .Z(n411) );
  GTECH_NOT U421 ( .A(I_a[2]), .Z(n239) );
  GTECH_AND_NOT U422 ( .A(I_b[2]), .B(n317), .Z(n416) );
  GTECH_NOT U423 ( .A(I_a[0]), .Z(n317) );
  GTECH_XOR2 U424 ( .A(n420), .B(n421), .Z(N141) );
  GTECH_AND_NOT U425 ( .A(I_a[1]), .B(n332), .Z(n421) );
  GTECH_NOT U426 ( .A(n422), .Z(n420) );
  GTECH_OR_NOT U427 ( .A(n258), .B(I_a[0]), .Z(n422) );
  GTECH_NOT U428 ( .A(I_b[1]), .Z(n258) );
  GTECH_AND_NOT U429 ( .A(I_a[0]), .B(n332), .Z(N140) );
  GTECH_NOT U430 ( .A(I_b[0]), .Z(n332) );
endmodule

