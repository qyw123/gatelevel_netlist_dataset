
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383;

  GTECH_MUX2 U138 ( .A(n277), .B(n278), .S(n279), .Z(sum[9]) );
  GTECH_XNOR2 U139 ( .A(n280), .B(n281), .Z(n278) );
  GTECH_XNOR2 U140 ( .A(n282), .B(n280), .Z(n277) );
  GTECH_OR_NOT U141 ( .A(n283), .B(n284), .Z(n280) );
  GTECH_NAND2 U142 ( .A(n285), .B(n286), .Z(sum[8]) );
  GTECH_OAI21 U143 ( .A(n282), .B(n287), .C(n279), .Z(n286) );
  GTECH_MUX2 U144 ( .A(n288), .B(n289), .S(n290), .Z(sum[7]) );
  GTECH_XNOR2 U145 ( .A(n291), .B(n292), .Z(n289) );
  GTECH_XOR2 U146 ( .A(n291), .B(n293), .Z(n288) );
  GTECH_AOI21 U147 ( .A(n294), .B(n295), .C(n296), .Z(n293) );
  GTECH_NOT U148 ( .A(n297), .Z(n296) );
  GTECH_XNOR2 U149 ( .A(a[7]), .B(b[7]), .Z(n291) );
  GTECH_MUX2 U150 ( .A(n298), .B(n299), .S(n300), .Z(sum[6]) );
  GTECH_XOR2 U151 ( .A(n295), .B(n301), .Z(n299) );
  GTECH_OAI21 U152 ( .A(n302), .B(n303), .C(n304), .Z(n295) );
  GTECH_XNOR2 U153 ( .A(n301), .B(n305), .Z(n298) );
  GTECH_AND2 U154 ( .A(n294), .B(n297), .Z(n301) );
  GTECH_MUX2 U155 ( .A(n306), .B(n307), .S(n308), .Z(sum[5]) );
  GTECH_OR_NOT U156 ( .A(n302), .B(n304), .Z(n308) );
  GTECH_OAI21 U157 ( .A(n309), .B(n300), .C(n303), .Z(n307) );
  GTECH_AO21 U158 ( .A(n303), .B(n300), .C(n309), .Z(n306) );
  GTECH_NOT U159 ( .A(n290), .Z(n300) );
  GTECH_XNOR2 U160 ( .A(n290), .B(n310), .Z(sum[4]) );
  GTECH_MUX2 U161 ( .A(n311), .B(n312), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U162 ( .A(n313), .B(n314), .Z(n312) );
  GTECH_XOR2 U163 ( .A(n313), .B(n315), .Z(n311) );
  GTECH_AOI21 U164 ( .A(n316), .B(n317), .C(n318), .Z(n315) );
  GTECH_NOT U165 ( .A(n319), .Z(n318) );
  GTECH_XNOR2 U166 ( .A(a[3]), .B(b[3]), .Z(n313) );
  GTECH_MUX2 U167 ( .A(n320), .B(n321), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U168 ( .A(n322), .B(n323), .Z(n321) );
  GTECH_XOR2 U169 ( .A(n317), .B(n322), .Z(n320) );
  GTECH_AND2 U170 ( .A(n316), .B(n319), .Z(n322) );
  GTECH_AO21 U171 ( .A(n324), .B(n325), .C(n326), .Z(n317) );
  GTECH_MUX2 U172 ( .A(n327), .B(n328), .S(n329), .Z(sum[1]) );
  GTECH_OR_NOT U173 ( .A(n326), .B(n324), .Z(n329) );
  GTECH_AO21 U174 ( .A(n330), .B(cin), .C(n325), .Z(n328) );
  GTECH_OAI21 U175 ( .A(cin), .B(n325), .C(n330), .Z(n327) );
  GTECH_AND2 U176 ( .A(b[0]), .B(a[0]), .Z(n325) );
  GTECH_MUX2 U177 ( .A(n331), .B(n332), .S(n333), .Z(sum[15]) );
  GTECH_XOR2 U178 ( .A(n334), .B(n335), .Z(n332) );
  GTECH_XOR2 U179 ( .A(n336), .B(n334), .Z(n331) );
  GTECH_XOR2 U180 ( .A(a[15]), .B(b[15]), .Z(n334) );
  GTECH_OA21 U181 ( .A(a[14]), .B(n337), .C(n338), .Z(n336) );
  GTECH_AO21 U182 ( .A(n337), .B(a[14]), .C(b[14]), .Z(n338) );
  GTECH_MUX2 U183 ( .A(n339), .B(n340), .S(n333), .Z(sum[14]) );
  GTECH_XOR2 U184 ( .A(n341), .B(n342), .Z(n340) );
  GTECH_XNOR2 U185 ( .A(n341), .B(n337), .Z(n339) );
  GTECH_AO21 U186 ( .A(n343), .B(n344), .C(n345), .Z(n337) );
  GTECH_XNOR2 U187 ( .A(n346), .B(n347), .Z(n341) );
  GTECH_MUX2 U188 ( .A(n348), .B(n349), .S(n333), .Z(sum[13]) );
  GTECH_XNOR2 U189 ( .A(n350), .B(n351), .Z(n349) );
  GTECH_XNOR2 U190 ( .A(n344), .B(n350), .Z(n348) );
  GTECH_OR_NOT U191 ( .A(n345), .B(n343), .Z(n350) );
  GTECH_NAND2 U192 ( .A(n352), .B(n353), .Z(sum[12]) );
  GTECH_OAI21 U193 ( .A(n344), .B(n354), .C(n333), .Z(n353) );
  GTECH_MUX2 U194 ( .A(n355), .B(n356), .S(n279), .Z(sum[11]) );
  GTECH_XNOR2 U195 ( .A(n357), .B(n358), .Z(n356) );
  GTECH_XOR2 U196 ( .A(n357), .B(n359), .Z(n355) );
  GTECH_AOI21 U197 ( .A(n360), .B(n361), .C(n362), .Z(n359) );
  GTECH_NOT U198 ( .A(n363), .Z(n362) );
  GTECH_XNOR2 U199 ( .A(a[11]), .B(b[11]), .Z(n357) );
  GTECH_MUX2 U200 ( .A(n364), .B(n365), .S(n279), .Z(sum[10]) );
  GTECH_XNOR2 U201 ( .A(n366), .B(n367), .Z(n365) );
  GTECH_XOR2 U202 ( .A(n361), .B(n366), .Z(n364) );
  GTECH_AND2 U203 ( .A(n360), .B(n363), .Z(n366) );
  GTECH_AO21 U204 ( .A(n284), .B(n282), .C(n283), .Z(n361) );
  GTECH_XOR2 U205 ( .A(cin), .B(n368), .Z(sum[0]) );
  GTECH_OAI21 U206 ( .A(n369), .B(n370), .C(n352), .Z(cout) );
  GTECH_OR3 U207 ( .A(n354), .B(n344), .C(n333), .Z(n352) );
  GTECH_NOT U208 ( .A(n369), .Z(n333) );
  GTECH_AND2 U209 ( .A(b[12]), .B(a[12]), .Z(n344) );
  GTECH_NOT U210 ( .A(n351), .Z(n354) );
  GTECH_AOI21 U211 ( .A(n335), .B(a[15]), .C(n371), .Z(n370) );
  GTECH_OA21 U212 ( .A(a[15]), .B(n335), .C(b[15]), .Z(n371) );
  GTECH_OAI21 U213 ( .A(n342), .B(n346), .C(n372), .Z(n335) );
  GTECH_AO21 U214 ( .A(n346), .B(n342), .C(n347), .Z(n372) );
  GTECH_NOT U215 ( .A(b[14]), .Z(n347) );
  GTECH_NOT U216 ( .A(a[14]), .Z(n346) );
  GTECH_AOI21 U217 ( .A(n351), .B(n343), .C(n345), .Z(n342) );
  GTECH_AND2 U218 ( .A(b[13]), .B(a[13]), .Z(n345) );
  GTECH_OR2 U219 ( .A(b[13]), .B(a[13]), .Z(n343) );
  GTECH_OR2 U220 ( .A(a[12]), .B(b[12]), .Z(n351) );
  GTECH_OA21 U221 ( .A(n373), .B(n374), .C(n285), .Z(n369) );
  GTECH_OR3 U222 ( .A(n287), .B(n282), .C(n279), .Z(n285) );
  GTECH_AND2 U223 ( .A(b[8]), .B(a[8]), .Z(n282) );
  GTECH_NOT U224 ( .A(n281), .Z(n287) );
  GTECH_NOT U225 ( .A(n279), .Z(n374) );
  GTECH_MUX2 U226 ( .A(n375), .B(n376), .S(n290), .Z(n279) );
  GTECH_MUX2 U227 ( .A(n368), .B(n377), .S(cin), .Z(n290) );
  GTECH_OA21 U228 ( .A(a[3]), .B(n314), .C(n378), .Z(n377) );
  GTECH_AO21 U229 ( .A(n314), .B(a[3]), .C(b[3]), .Z(n378) );
  GTECH_OAI21 U230 ( .A(n323), .B(n379), .C(n319), .Z(n314) );
  GTECH_NAND2 U231 ( .A(b[2]), .B(a[2]), .Z(n319) );
  GTECH_NOT U232 ( .A(n316), .Z(n379) );
  GTECH_OR2 U233 ( .A(b[2]), .B(a[2]), .Z(n316) );
  GTECH_AOI21 U234 ( .A(n324), .B(n330), .C(n326), .Z(n323) );
  GTECH_AND2 U235 ( .A(a[1]), .B(b[1]), .Z(n326) );
  GTECH_OR2 U236 ( .A(b[0]), .B(a[0]), .Z(n330) );
  GTECH_OR2 U237 ( .A(a[1]), .B(b[1]), .Z(n324) );
  GTECH_XOR2 U238 ( .A(a[0]), .B(b[0]), .Z(n368) );
  GTECH_OA21 U239 ( .A(a[7]), .B(n292), .C(n380), .Z(n376) );
  GTECH_AO21 U240 ( .A(n292), .B(a[7]), .C(b[7]), .Z(n380) );
  GTECH_OAI21 U241 ( .A(n305), .B(n381), .C(n297), .Z(n292) );
  GTECH_NAND2 U242 ( .A(a[6]), .B(b[6]), .Z(n297) );
  GTECH_NOT U243 ( .A(n294), .Z(n381) );
  GTECH_OR2 U244 ( .A(b[6]), .B(a[6]), .Z(n294) );
  GTECH_OA21 U245 ( .A(n302), .B(n309), .C(n304), .Z(n305) );
  GTECH_NAND2 U246 ( .A(b[5]), .B(a[5]), .Z(n304) );
  GTECH_NOR2 U247 ( .A(a[5]), .B(b[5]), .Z(n302) );
  GTECH_NOT U248 ( .A(n310), .Z(n375) );
  GTECH_OR_NOT U249 ( .A(n309), .B(n303), .Z(n310) );
  GTECH_NAND2 U250 ( .A(b[4]), .B(a[4]), .Z(n303) );
  GTECH_NOR2 U251 ( .A(a[4]), .B(b[4]), .Z(n309) );
  GTECH_AOI21 U252 ( .A(n358), .B(a[11]), .C(n382), .Z(n373) );
  GTECH_OA21 U253 ( .A(a[11]), .B(n358), .C(b[11]), .Z(n382) );
  GTECH_OAI21 U254 ( .A(n367), .B(n383), .C(n363), .Z(n358) );
  GTECH_NAND2 U255 ( .A(a[10]), .B(b[10]), .Z(n363) );
  GTECH_NOT U256 ( .A(n360), .Z(n383) );
  GTECH_OR2 U257 ( .A(b[10]), .B(a[10]), .Z(n360) );
  GTECH_AOI21 U258 ( .A(n284), .B(n281), .C(n283), .Z(n367) );
  GTECH_AND2 U259 ( .A(b[9]), .B(a[9]), .Z(n283) );
  GTECH_OR2 U260 ( .A(a[8]), .B(b[8]), .Z(n281) );
  GTECH_OR2 U261 ( .A(a[9]), .B(b[9]), .Z(n284) );
endmodule

