
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387;

  GTECH_MUX2 U132 ( .A(n271), .B(n272), .S(n273), .Z(sum[9]) );
  GTECH_XNOR2 U133 ( .A(n274), .B(n275), .Z(n272) );
  GTECH_XOR2 U134 ( .A(n275), .B(n276), .Z(n271) );
  GTECH_OA21 U135 ( .A(b[9]), .B(a[9]), .C(n277), .Z(n275) );
  GTECH_NAND2 U136 ( .A(n278), .B(n279), .Z(sum[8]) );
  GTECH_OAI21 U137 ( .A(n280), .B(n281), .C(n282), .Z(n279) );
  GTECH_MUX2 U138 ( .A(n283), .B(n284), .S(n285), .Z(sum[7]) );
  GTECH_XNOR2 U139 ( .A(n286), .B(n287), .Z(n284) );
  GTECH_XOR2 U140 ( .A(n286), .B(n288), .Z(n283) );
  GTECH_OA21 U141 ( .A(n289), .B(n290), .C(n291), .Z(n288) );
  GTECH_ADD_AB U142 ( .A(n292), .B(n293), .COUT(n289) );
  GTECH_XNOR2 U143 ( .A(a[7]), .B(b[7]), .Z(n286) );
  GTECH_MUX2 U144 ( .A(n294), .B(n295), .S(n285), .Z(sum[6]) );
  GTECH_XOR2 U145 ( .A(n296), .B(n297), .Z(n295) );
  GTECH_XOR2 U146 ( .A(n296), .B(n290), .Z(n294) );
  GTECH_ADD_AB U147 ( .A(n298), .B(n299), .COUT(n290) );
  GTECH_OAI21 U148 ( .A(b[5]), .B(a[5]), .C(n300), .Z(n299) );
  GTECH_OAI21 U149 ( .A(b[6]), .B(a[6]), .C(n291), .Z(n296) );
  GTECH_NOT U150 ( .A(n301), .Z(n291) );
  GTECH_MUX2 U151 ( .A(n302), .B(n303), .S(n304), .Z(sum[5]) );
  GTECH_OA21 U152 ( .A(b[5]), .B(a[5]), .C(n298), .Z(n304) );
  GTECH_OAI21 U153 ( .A(n300), .B(n285), .C(n305), .Z(n303) );
  GTECH_AO21 U154 ( .A(n305), .B(n285), .C(n300), .Z(n302) );
  GTECH_XNOR2 U155 ( .A(n285), .B(n306), .Z(sum[4]) );
  GTECH_MUX2 U156 ( .A(n307), .B(n308), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U157 ( .A(n309), .B(n310), .Z(n308) );
  GTECH_XOR2 U158 ( .A(n309), .B(n311), .Z(n307) );
  GTECH_OA21 U159 ( .A(n312), .B(n313), .C(n314), .Z(n311) );
  GTECH_ADD_AB U160 ( .A(n315), .B(n316), .COUT(n312) );
  GTECH_XNOR2 U161 ( .A(a[3]), .B(b[3]), .Z(n309) );
  GTECH_MUX2 U162 ( .A(n317), .B(n318), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U163 ( .A(n319), .B(n320), .Z(n318) );
  GTECH_XOR2 U164 ( .A(n319), .B(n313), .Z(n317) );
  GTECH_ADD_AB U165 ( .A(n321), .B(n322), .COUT(n313) );
  GTECH_OAI21 U166 ( .A(b[1]), .B(a[1]), .C(n323), .Z(n322) );
  GTECH_OAI21 U167 ( .A(b[2]), .B(a[2]), .C(n314), .Z(n319) );
  GTECH_NOT U168 ( .A(n324), .Z(n314) );
  GTECH_MUX2 U169 ( .A(n325), .B(n326), .S(n327), .Z(sum[1]) );
  GTECH_OA21 U170 ( .A(b[1]), .B(a[1]), .C(n321), .Z(n327) );
  GTECH_OAI21 U171 ( .A(cin), .B(n323), .C(n328), .Z(n326) );
  GTECH_AO21 U172 ( .A(n328), .B(cin), .C(n323), .Z(n325) );
  GTECH_ADD_AB U173 ( .A(a[0]), .B(b[0]), .COUT(n323) );
  GTECH_MUX2 U174 ( .A(n329), .B(n330), .S(n331), .Z(sum[15]) );
  GTECH_XOR2 U175 ( .A(n332), .B(n333), .Z(n330) );
  GTECH_OA21 U176 ( .A(n334), .B(n335), .C(n336), .Z(n333) );
  GTECH_NOR2 U177 ( .A(a[14]), .B(b[14]), .Z(n334) );
  GTECH_XNOR2 U178 ( .A(n332), .B(n337), .Z(n329) );
  GTECH_XNOR2 U179 ( .A(a[15]), .B(b[15]), .Z(n332) );
  GTECH_MUX2 U180 ( .A(n338), .B(n339), .S(n331), .Z(sum[14]) );
  GTECH_XOR2 U181 ( .A(n340), .B(n335), .Z(n339) );
  GTECH_ADD_AB U182 ( .A(n341), .B(n342), .COUT(n335) );
  GTECH_OAI21 U183 ( .A(b[13]), .B(a[13]), .C(n343), .Z(n342) );
  GTECH_XNOR2 U184 ( .A(n340), .B(n344), .Z(n338) );
  GTECH_OAI21 U185 ( .A(b[14]), .B(a[14]), .C(n336), .Z(n340) );
  GTECH_MUX2 U186 ( .A(n345), .B(n346), .S(n331), .Z(sum[13]) );
  GTECH_XOR2 U187 ( .A(n347), .B(n348), .Z(n346) );
  GTECH_XNOR2 U188 ( .A(n348), .B(n349), .Z(n345) );
  GTECH_OAI21 U189 ( .A(b[13]), .B(a[13]), .C(n341), .Z(n348) );
  GTECH_NAND2 U190 ( .A(n350), .B(n351), .Z(sum[12]) );
  GTECH_OAI21 U191 ( .A(n343), .B(n352), .C(n353), .Z(n351) );
  GTECH_MUX2 U192 ( .A(n354), .B(n355), .S(n273), .Z(sum[11]) );
  GTECH_XOR2 U193 ( .A(n356), .B(n357), .Z(n355) );
  GTECH_OA21 U194 ( .A(n358), .B(n359), .C(n360), .Z(n357) );
  GTECH_ADD_AB U195 ( .A(n361), .B(n362), .COUT(n358) );
  GTECH_XNOR2 U196 ( .A(n356), .B(n363), .Z(n354) );
  GTECH_XNOR2 U197 ( .A(a[11]), .B(b[11]), .Z(n356) );
  GTECH_MUX2 U198 ( .A(n364), .B(n365), .S(n273), .Z(sum[10]) );
  GTECH_XOR2 U199 ( .A(n366), .B(n359), .Z(n365) );
  GTECH_ADD_AB U200 ( .A(n277), .B(n367), .COUT(n359) );
  GTECH_OAI21 U201 ( .A(b[9]), .B(a[9]), .C(n280), .Z(n367) );
  GTECH_XOR2 U202 ( .A(n366), .B(n368), .Z(n364) );
  GTECH_OAI21 U203 ( .A(b[10]), .B(a[10]), .C(n360), .Z(n366) );
  GTECH_NOT U204 ( .A(n369), .Z(n360) );
  GTECH_XOR2 U205 ( .A(cin), .B(n370), .Z(sum[0]) );
  GTECH_OAI21 U206 ( .A(n331), .B(n371), .C(n350), .Z(cout) );
  GTECH_NAND3 U207 ( .A(n347), .B(n349), .C(n331), .Z(n350) );
  GTECH_NOT U208 ( .A(n343), .Z(n347) );
  GTECH_ADD_AB U209 ( .A(b[12]), .B(a[12]), .COUT(n343) );
  GTECH_AOI21 U210 ( .A(n337), .B(a[15]), .C(n372), .Z(n371) );
  GTECH_OA21 U211 ( .A(a[15]), .B(n337), .C(b[15]), .Z(n372) );
  GTECH_NAND2 U212 ( .A(n336), .B(n373), .Z(n337) );
  GTECH_OAI21 U213 ( .A(a[14]), .B(b[14]), .C(n344), .Z(n373) );
  GTECH_NAND2 U214 ( .A(n341), .B(n374), .Z(n344) );
  GTECH_OAI21 U215 ( .A(a[13]), .B(b[13]), .C(n349), .Z(n374) );
  GTECH_NOT U216 ( .A(n352), .Z(n349) );
  GTECH_NOR2 U217 ( .A(a[12]), .B(b[12]), .Z(n352) );
  GTECH_NAND2 U218 ( .A(b[13]), .B(a[13]), .Z(n341) );
  GTECH_NAND2 U219 ( .A(b[14]), .B(a[14]), .Z(n336) );
  GTECH_NOT U220 ( .A(n353), .Z(n331) );
  GTECH_OAI21 U221 ( .A(n375), .B(n273), .C(n278), .Z(n353) );
  GTECH_NAND3 U222 ( .A(n274), .B(n276), .C(n273), .Z(n278) );
  GTECH_NOT U223 ( .A(n280), .Z(n274) );
  GTECH_ADD_AB U224 ( .A(b[8]), .B(a[8]), .COUT(n280) );
  GTECH_NOT U225 ( .A(n282), .Z(n273) );
  GTECH_MUX2 U226 ( .A(n376), .B(n377), .S(n285), .Z(n282) );
  GTECH_MUX2 U227 ( .A(n370), .B(n378), .S(cin), .Z(n285) );
  GTECH_OA21 U228 ( .A(a[3]), .B(n310), .C(n379), .Z(n378) );
  GTECH_AO21 U229 ( .A(n310), .B(a[3]), .C(b[3]), .Z(n379) );
  GTECH_OR_NOT U230 ( .A(n324), .B(n380), .Z(n310) );
  GTECH_AO21 U231 ( .A(n315), .B(n316), .C(n320), .Z(n380) );
  GTECH_ADD_AB U232 ( .A(n321), .B(n381), .COUT(n320) );
  GTECH_OAI21 U233 ( .A(a[1]), .B(b[1]), .C(n328), .Z(n381) );
  GTECH_OR2 U234 ( .A(b[0]), .B(a[0]), .Z(n328) );
  GTECH_NAND2 U235 ( .A(b[1]), .B(a[1]), .Z(n321) );
  GTECH_NOT U236 ( .A(b[2]), .Z(n316) );
  GTECH_NOT U237 ( .A(a[2]), .Z(n315) );
  GTECH_ADD_AB U238 ( .A(b[2]), .B(a[2]), .COUT(n324) );
  GTECH_XOR2 U239 ( .A(a[0]), .B(b[0]), .Z(n370) );
  GTECH_OA21 U240 ( .A(a[7]), .B(n287), .C(n382), .Z(n377) );
  GTECH_AO21 U241 ( .A(n287), .B(a[7]), .C(b[7]), .Z(n382) );
  GTECH_OR_NOT U242 ( .A(n301), .B(n383), .Z(n287) );
  GTECH_AO21 U243 ( .A(n292), .B(n293), .C(n297), .Z(n383) );
  GTECH_ADD_AB U244 ( .A(n298), .B(n384), .COUT(n297) );
  GTECH_OAI21 U245 ( .A(a[5]), .B(b[5]), .C(n305), .Z(n384) );
  GTECH_NAND2 U246 ( .A(b[5]), .B(a[5]), .Z(n298) );
  GTECH_NOT U247 ( .A(b[6]), .Z(n293) );
  GTECH_NOT U248 ( .A(a[6]), .Z(n292) );
  GTECH_ADD_AB U249 ( .A(b[6]), .B(a[6]), .COUT(n301) );
  GTECH_NOT U250 ( .A(n306), .Z(n376) );
  GTECH_OR_NOT U251 ( .A(n300), .B(n305), .Z(n306) );
  GTECH_OR2 U252 ( .A(a[4]), .B(b[4]), .Z(n305) );
  GTECH_ADD_AB U253 ( .A(b[4]), .B(a[4]), .COUT(n300) );
  GTECH_AOI21 U254 ( .A(n363), .B(a[11]), .C(n385), .Z(n375) );
  GTECH_OA21 U255 ( .A(a[11]), .B(n363), .C(b[11]), .Z(n385) );
  GTECH_OR_NOT U256 ( .A(n369), .B(n386), .Z(n363) );
  GTECH_AO21 U257 ( .A(n361), .B(n362), .C(n368), .Z(n386) );
  GTECH_ADD_AB U258 ( .A(n277), .B(n387), .COUT(n368) );
  GTECH_OAI21 U259 ( .A(a[9]), .B(b[9]), .C(n276), .Z(n387) );
  GTECH_NOT U260 ( .A(n281), .Z(n276) );
  GTECH_NOR2 U261 ( .A(a[8]), .B(b[8]), .Z(n281) );
  GTECH_NAND2 U262 ( .A(b[9]), .B(a[9]), .Z(n277) );
  GTECH_NOT U263 ( .A(b[10]), .Z(n362) );
  GTECH_NOT U264 ( .A(a[10]), .Z(n361) );
  GTECH_ADD_AB U265 ( .A(b[10]), .B(a[10]), .COUT(n369) );
endmodule

