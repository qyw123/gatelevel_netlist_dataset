
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NAND2 U83 ( .A(n93), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI21 U86 ( .A(n98), .B(n99), .C(n100), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_NOT U88 ( .A(n102), .Z(n98) );
  GTECH_NAND2 U89 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n104), .Z(n84) );
  GTECH_NAND2 U91 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_XOR2 U92 ( .A(n106), .B(n105), .Z(N153) );
  GTECH_NOT U93 ( .A(n107), .Z(n105) );
  GTECH_XOR3 U94 ( .A(n108), .B(n93), .C(n95), .Z(n107) );
  GTECH_XOR3 U95 ( .A(n101), .B(n103), .C(n102), .Z(n95) );
  GTECH_OAI21 U96 ( .A(n109), .B(n110), .C(n111), .Z(n102) );
  GTECH_OAI21 U97 ( .A(n112), .B(n113), .C(n114), .Z(n111) );
  GTECH_NOT U98 ( .A(n113), .Z(n109) );
  GTECH_NOT U99 ( .A(n115), .Z(n103) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n115) );
  GTECH_NOT U101 ( .A(n99), .Z(n101) );
  GTECH_NAND2 U102 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U103 ( .A(n116), .B(n117), .C(n118), .COUT(n93) );
  GTECH_NOT U104 ( .A(n119), .Z(n118) );
  GTECH_XOR2 U105 ( .A(n120), .B(n121), .Z(n117) );
  GTECH_AND2 U106 ( .A(I_a[7]), .B(I_b[5]), .Z(n121) );
  GTECH_NOT U107 ( .A(n122), .Z(n120) );
  GTECH_NOT U108 ( .A(n94), .Z(n108) );
  GTECH_NAND2 U109 ( .A(I_a[7]), .B(n122), .Z(n94) );
  GTECH_NOT U110 ( .A(n123), .Z(n106) );
  GTECH_NAND2 U111 ( .A(n124), .B(n125), .Z(n123) );
  GTECH_NOT U112 ( .A(n126), .Z(n125) );
  GTECH_XOR2 U113 ( .A(n126), .B(n127), .Z(N152) );
  GTECH_NOT U114 ( .A(n124), .Z(n127) );
  GTECH_XNOR4 U115 ( .A(n128), .B(n119), .C(n122), .D(n116), .Z(n124) );
  GTECH_ADD_ABC U116 ( .A(n129), .B(n130), .C(n131), .COUT(n116) );
  GTECH_NOT U117 ( .A(n132), .Z(n131) );
  GTECH_XOR3 U118 ( .A(n133), .B(n134), .C(n135), .Z(n130) );
  GTECH_OAI21 U119 ( .A(n135), .B(n136), .C(n137), .Z(n122) );
  GTECH_OAI21 U120 ( .A(n133), .B(n138), .C(n134), .Z(n137) );
  GTECH_NOT U121 ( .A(n138), .Z(n135) );
  GTECH_XOR3 U122 ( .A(n112), .B(n114), .C(n113), .Z(n119) );
  GTECH_OAI21 U123 ( .A(n139), .B(n140), .C(n141), .Z(n113) );
  GTECH_OAI21 U124 ( .A(n142), .B(n143), .C(n144), .Z(n141) );
  GTECH_NOT U125 ( .A(n143), .Z(n139) );
  GTECH_NOT U126 ( .A(n145), .Z(n114) );
  GTECH_NAND2 U127 ( .A(I_b[7]), .B(I_a[5]), .Z(n145) );
  GTECH_NOT U128 ( .A(n110), .Z(n112) );
  GTECH_NAND2 U129 ( .A(I_b[6]), .B(I_a[6]), .Z(n110) );
  GTECH_AND2 U130 ( .A(I_a[7]), .B(I_b[5]), .Z(n128) );
  GTECH_ADD_ABC U131 ( .A(n146), .B(n147), .C(n148), .COUT(n126) );
  GTECH_NOT U132 ( .A(n149), .Z(n148) );
  GTECH_OA22 U133 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n147) );
  GTECH_OA22 U134 ( .A(n154), .B(n155), .C(n156), .D(n157), .Z(n146) );
  GTECH_AND2 U135 ( .A(n156), .B(n157), .Z(n154) );
  GTECH_XOR3 U136 ( .A(n158), .B(n149), .C(n159), .Z(N151) );
  GTECH_AOI2N2 U137 ( .A(n160), .B(n161), .C(n156), .D(n157), .Z(n159) );
  GTECH_OR_NOT U138 ( .A(n162), .B(n157), .Z(n161) );
  GTECH_XOR2 U139 ( .A(n163), .B(n129), .Z(n149) );
  GTECH_ADD_ABC U140 ( .A(n164), .B(n165), .C(n166), .COUT(n129) );
  GTECH_NOT U141 ( .A(n167), .Z(n166) );
  GTECH_XOR3 U142 ( .A(n168), .B(n169), .C(n170), .Z(n165) );
  GTECH_XNOR4 U143 ( .A(n134), .B(n138), .C(n132), .D(n133), .Z(n163) );
  GTECH_NOT U144 ( .A(n136), .Z(n133) );
  GTECH_NAND2 U145 ( .A(I_a[7]), .B(I_b[4]), .Z(n136) );
  GTECH_XOR3 U146 ( .A(n142), .B(n144), .C(n143), .Z(n132) );
  GTECH_OAI21 U147 ( .A(n171), .B(n172), .C(n173), .Z(n143) );
  GTECH_OAI21 U148 ( .A(n174), .B(n175), .C(n176), .Z(n173) );
  GTECH_NOT U149 ( .A(n175), .Z(n171) );
  GTECH_NOT U150 ( .A(n177), .Z(n144) );
  GTECH_NAND2 U151 ( .A(I_b[7]), .B(I_a[4]), .Z(n177) );
  GTECH_NOT U152 ( .A(n140), .Z(n142) );
  GTECH_NAND2 U153 ( .A(I_b[6]), .B(I_a[5]), .Z(n140) );
  GTECH_OAI21 U154 ( .A(n170), .B(n178), .C(n179), .Z(n138) );
  GTECH_OAI21 U155 ( .A(n168), .B(n180), .C(n169), .Z(n179) );
  GTECH_NOT U156 ( .A(n180), .Z(n170) );
  GTECH_NOT U157 ( .A(n181), .Z(n134) );
  GTECH_NAND2 U158 ( .A(I_a[6]), .B(I_b[5]), .Z(n181) );
  GTECH_OA22 U159 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n158) );
  GTECH_NOT U160 ( .A(n182), .Z(n153) );
  GTECH_NOT U161 ( .A(I_a[7]), .Z(n151) );
  GTECH_XOR3 U162 ( .A(n156), .B(n183), .C(n155), .Z(N150) );
  GTECH_NOT U163 ( .A(n160), .Z(n155) );
  GTECH_XOR2 U164 ( .A(n184), .B(n164), .Z(n160) );
  GTECH_ADD_ABC U165 ( .A(n185), .B(n186), .C(n187), .COUT(n164) );
  GTECH_NOT U166 ( .A(n188), .Z(n187) );
  GTECH_XOR3 U167 ( .A(n189), .B(n190), .C(n191), .Z(n186) );
  GTECH_XNOR4 U168 ( .A(n169), .B(n180), .C(n167), .D(n168), .Z(n184) );
  GTECH_NOT U169 ( .A(n178), .Z(n168) );
  GTECH_NAND2 U170 ( .A(I_a[6]), .B(I_b[4]), .Z(n178) );
  GTECH_XOR3 U171 ( .A(n174), .B(n176), .C(n175), .Z(n167) );
  GTECH_OAI21 U172 ( .A(n192), .B(n193), .C(n194), .Z(n175) );
  GTECH_OAI21 U173 ( .A(n195), .B(n196), .C(n197), .Z(n194) );
  GTECH_NOT U174 ( .A(n196), .Z(n192) );
  GTECH_NOT U175 ( .A(n198), .Z(n176) );
  GTECH_NAND2 U176 ( .A(I_b[7]), .B(I_a[3]), .Z(n198) );
  GTECH_NOT U177 ( .A(n172), .Z(n174) );
  GTECH_NAND2 U178 ( .A(I_b[6]), .B(I_a[4]), .Z(n172) );
  GTECH_OAI21 U179 ( .A(n191), .B(n199), .C(n200), .Z(n180) );
  GTECH_OAI21 U180 ( .A(n189), .B(n201), .C(n190), .Z(n200) );
  GTECH_NOT U181 ( .A(n201), .Z(n191) );
  GTECH_NOT U182 ( .A(n202), .Z(n169) );
  GTECH_NAND2 U183 ( .A(I_a[5]), .B(I_b[5]), .Z(n202) );
  GTECH_NOT U184 ( .A(n157), .Z(n183) );
  GTECH_XOR2 U185 ( .A(n182), .B(n152), .Z(n157) );
  GTECH_AOI2N2 U186 ( .A(n203), .B(n204), .C(n205), .D(n206), .Z(n152) );
  GTECH_NAND2 U187 ( .A(n205), .B(n206), .Z(n204) );
  GTECH_XOR2 U188 ( .A(n207), .B(n150), .Z(n182) );
  GTECH_AND2 U189 ( .A(n208), .B(n209), .Z(n150) );
  GTECH_OR_NOT U190 ( .A(n210), .B(n211), .Z(n209) );
  GTECH_OAI21 U191 ( .A(n212), .B(n211), .C(n213), .Z(n208) );
  GTECH_NAND2 U192 ( .A(I_a[7]), .B(I_b[3]), .Z(n207) );
  GTECH_NOT U193 ( .A(n162), .Z(n156) );
  GTECH_OAI2N2 U194 ( .A(n214), .B(n215), .C(n216), .D(n217), .Z(n162) );
  GTECH_NAND2 U195 ( .A(n214), .B(n215), .Z(n217) );
  GTECH_XOR3 U196 ( .A(n214), .B(n218), .C(n219), .Z(N149) );
  GTECH_NOT U197 ( .A(n216), .Z(n219) );
  GTECH_XOR2 U198 ( .A(n220), .B(n185), .Z(n216) );
  GTECH_ADD_ABC U199 ( .A(n221), .B(n222), .C(n223), .COUT(n185) );
  GTECH_XOR3 U200 ( .A(n224), .B(n225), .C(n226), .Z(n222) );
  GTECH_OA22 U201 ( .A(n227), .B(n228), .C(n229), .D(n230), .Z(n221) );
  GTECH_AND2 U202 ( .A(n229), .B(n230), .Z(n227) );
  GTECH_XNOR4 U203 ( .A(n190), .B(n201), .C(n188), .D(n189), .Z(n220) );
  GTECH_NOT U204 ( .A(n199), .Z(n189) );
  GTECH_NAND2 U205 ( .A(I_a[5]), .B(I_b[4]), .Z(n199) );
  GTECH_XOR3 U206 ( .A(n195), .B(n197), .C(n196), .Z(n188) );
  GTECH_OAI21 U207 ( .A(n231), .B(n232), .C(n233), .Z(n196) );
  GTECH_NOT U208 ( .A(n234), .Z(n197) );
  GTECH_NAND2 U209 ( .A(I_b[7]), .B(I_a[2]), .Z(n234) );
  GTECH_NOT U210 ( .A(n193), .Z(n195) );
  GTECH_NAND2 U211 ( .A(I_b[6]), .B(I_a[3]), .Z(n193) );
  GTECH_OAI21 U212 ( .A(n226), .B(n235), .C(n236), .Z(n201) );
  GTECH_OAI21 U213 ( .A(n224), .B(n237), .C(n225), .Z(n236) );
  GTECH_NOT U214 ( .A(n237), .Z(n226) );
  GTECH_NOT U215 ( .A(n238), .Z(n190) );
  GTECH_NAND2 U216 ( .A(I_b[5]), .B(I_a[4]), .Z(n238) );
  GTECH_NOT U217 ( .A(n215), .Z(n218) );
  GTECH_XOR3 U218 ( .A(n239), .B(n205), .C(n203), .Z(n215) );
  GTECH_XOR3 U219 ( .A(n212), .B(n213), .C(n211), .Z(n203) );
  GTECH_OAI21 U220 ( .A(n240), .B(n241), .C(n242), .Z(n211) );
  GTECH_OAI21 U221 ( .A(n243), .B(n244), .C(n245), .Z(n242) );
  GTECH_NOT U222 ( .A(n244), .Z(n240) );
  GTECH_NOT U223 ( .A(n246), .Z(n213) );
  GTECH_NAND2 U224 ( .A(I_a[6]), .B(I_b[3]), .Z(n246) );
  GTECH_NOT U225 ( .A(n210), .Z(n212) );
  GTECH_NAND2 U226 ( .A(I_a[7]), .B(I_b[2]), .Z(n210) );
  GTECH_ADD_ABC U227 ( .A(n247), .B(n248), .C(n249), .COUT(n205) );
  GTECH_XOR2 U228 ( .A(n250), .B(n251), .Z(n248) );
  GTECH_AND2 U229 ( .A(I_a[7]), .B(I_b[1]), .Z(n251) );
  GTECH_NOT U230 ( .A(n206), .Z(n239) );
  GTECH_NAND2 U231 ( .A(I_a[7]), .B(n252), .Z(n206) );
  GTECH_ADD_ABC U232 ( .A(n253), .B(n254), .C(n255), .COUT(n214) );
  GTECH_XOR3 U233 ( .A(n247), .B(n256), .C(n249), .Z(n254) );
  GTECH_NOT U234 ( .A(n257), .Z(n249) );
  GTECH_XOR3 U235 ( .A(n258), .B(n255), .C(n253), .Z(N148) );
  GTECH_ADD_ABC U236 ( .A(n259), .B(n260), .C(n261), .COUT(n253) );
  GTECH_NOT U237 ( .A(n262), .Z(n261) );
  GTECH_XOR3 U238 ( .A(n263), .B(n264), .C(n265), .Z(n260) );
  GTECH_XOR2 U239 ( .A(n266), .B(n267), .Z(n255) );
  GTECH_OA22 U240 ( .A(n229), .B(n230), .C(n268), .D(n228), .Z(n267) );
  GTECH_AND_NOT U241 ( .A(n229), .B(n269), .Z(n268) );
  GTECH_XNOR4 U242 ( .A(n225), .B(n237), .C(n223), .D(n224), .Z(n266) );
  GTECH_NOT U243 ( .A(n235), .Z(n224) );
  GTECH_NAND2 U244 ( .A(I_b[4]), .B(I_a[4]), .Z(n235) );
  GTECH_XOR3 U245 ( .A(n270), .B(n271), .C(n233), .Z(n223) );
  GTECH_NAND3 U246 ( .A(I_b[6]), .B(I_a[1]), .C(n272), .Z(n233) );
  GTECH_NOT U247 ( .A(n232), .Z(n271) );
  GTECH_NAND2 U248 ( .A(I_b[7]), .B(I_a[1]), .Z(n232) );
  GTECH_NOT U249 ( .A(n231), .Z(n270) );
  GTECH_NAND2 U250 ( .A(I_b[6]), .B(I_a[2]), .Z(n231) );
  GTECH_OAI21 U251 ( .A(n273), .B(n274), .C(n275), .Z(n237) );
  GTECH_OAI21 U252 ( .A(n276), .B(n277), .C(n278), .Z(n275) );
  GTECH_NOT U253 ( .A(n277), .Z(n273) );
  GTECH_NOT U254 ( .A(n279), .Z(n225) );
  GTECH_NAND2 U255 ( .A(I_b[5]), .B(I_a[3]), .Z(n279) );
  GTECH_XOR3 U256 ( .A(n256), .B(n257), .C(n247), .Z(n258) );
  GTECH_ADD_ABC U257 ( .A(n263), .B(n280), .C(n265), .COUT(n247) );
  GTECH_NOT U258 ( .A(n281), .Z(n265) );
  GTECH_XOR3 U259 ( .A(n282), .B(n283), .C(n284), .Z(n280) );
  GTECH_XOR3 U260 ( .A(n243), .B(n245), .C(n244), .Z(n257) );
  GTECH_OAI21 U261 ( .A(n285), .B(n286), .C(n287), .Z(n244) );
  GTECH_OAI21 U262 ( .A(n288), .B(n289), .C(n290), .Z(n287) );
  GTECH_NOT U263 ( .A(n289), .Z(n285) );
  GTECH_NOT U264 ( .A(n291), .Z(n245) );
  GTECH_NAND2 U265 ( .A(I_a[5]), .B(I_b[3]), .Z(n291) );
  GTECH_NOT U266 ( .A(n241), .Z(n243) );
  GTECH_NAND2 U267 ( .A(I_a[6]), .B(I_b[2]), .Z(n241) );
  GTECH_XOR2 U268 ( .A(n292), .B(n250), .Z(n256) );
  GTECH_NOT U269 ( .A(n252), .Z(n250) );
  GTECH_OAI21 U270 ( .A(n284), .B(n293), .C(n294), .Z(n252) );
  GTECH_OAI21 U271 ( .A(n282), .B(n295), .C(n283), .Z(n294) );
  GTECH_NOT U272 ( .A(n295), .Z(n284) );
  GTECH_AND2 U273 ( .A(I_a[7]), .B(I_b[1]), .Z(n292) );
  GTECH_XOR2 U274 ( .A(n296), .B(n259), .Z(N147) );
  GTECH_ADD_ABC U275 ( .A(n297), .B(n298), .C(n299), .COUT(n259) );
  GTECH_XOR3 U276 ( .A(n300), .B(n301), .C(n302), .Z(n298) );
  GTECH_NOT U277 ( .A(n303), .Z(n301) );
  GTECH_OA22 U278 ( .A(n304), .B(n305), .C(n306), .D(n307), .Z(n297) );
  GTECH_AND2 U279 ( .A(n306), .B(n307), .Z(n304) );
  GTECH_XNOR4 U280 ( .A(n264), .B(n281), .C(n262), .D(n263), .Z(n296) );
  GTECH_ADD_ABC U281 ( .A(n300), .B(n308), .C(n302), .COUT(n263) );
  GTECH_NOT U282 ( .A(n309), .Z(n302) );
  GTECH_XOR3 U283 ( .A(n310), .B(n311), .C(n312), .Z(n308) );
  GTECH_XOR3 U284 ( .A(n313), .B(n230), .C(n229), .Z(n262) );
  GTECH_XOR2 U285 ( .A(n314), .B(n272), .Z(n229) );
  GTECH_NOT U286 ( .A(n315), .Z(n272) );
  GTECH_NAND2 U287 ( .A(I_b[7]), .B(I_a[0]), .Z(n315) );
  GTECH_NAND2 U288 ( .A(I_b[6]), .B(I_a[1]), .Z(n314) );
  GTECH_NOT U289 ( .A(n269), .Z(n230) );
  GTECH_XOR3 U290 ( .A(n276), .B(n278), .C(n277), .Z(n269) );
  GTECH_OAI21 U291 ( .A(n316), .B(n317), .C(n318), .Z(n277) );
  GTECH_NOT U292 ( .A(n319), .Z(n278) );
  GTECH_NAND2 U293 ( .A(I_b[5]), .B(I_a[2]), .Z(n319) );
  GTECH_NOT U294 ( .A(n274), .Z(n276) );
  GTECH_NAND2 U295 ( .A(I_b[4]), .B(I_a[3]), .Z(n274) );
  GTECH_NOT U296 ( .A(n228), .Z(n313) );
  GTECH_NAND3 U297 ( .A(I_a[0]), .B(n320), .C(I_b[6]), .Z(n228) );
  GTECH_NOT U298 ( .A(n321), .Z(n320) );
  GTECH_XOR3 U299 ( .A(n288), .B(n290), .C(n289), .Z(n281) );
  GTECH_OAI21 U300 ( .A(n322), .B(n323), .C(n324), .Z(n289) );
  GTECH_OAI21 U301 ( .A(n325), .B(n326), .C(n327), .Z(n324) );
  GTECH_NOT U302 ( .A(n326), .Z(n322) );
  GTECH_NOT U303 ( .A(n328), .Z(n290) );
  GTECH_NAND2 U304 ( .A(I_b[3]), .B(I_a[4]), .Z(n328) );
  GTECH_NOT U305 ( .A(n286), .Z(n288) );
  GTECH_NAND2 U306 ( .A(I_a[5]), .B(I_b[2]), .Z(n286) );
  GTECH_NOT U307 ( .A(n329), .Z(n264) );
  GTECH_XOR3 U308 ( .A(n282), .B(n283), .C(n295), .Z(n329) );
  GTECH_OAI21 U309 ( .A(n312), .B(n330), .C(n331), .Z(n295) );
  GTECH_OAI21 U310 ( .A(n310), .B(n332), .C(n311), .Z(n331) );
  GTECH_NOT U311 ( .A(n332), .Z(n312) );
  GTECH_NOT U312 ( .A(n333), .Z(n283) );
  GTECH_NAND2 U313 ( .A(I_a[6]), .B(I_b[1]), .Z(n333) );
  GTECH_NOT U314 ( .A(n293), .Z(n282) );
  GTECH_NAND2 U315 ( .A(I_a[7]), .B(I_b[0]), .Z(n293) );
  GTECH_XOR2 U316 ( .A(n334), .B(n335), .Z(N146) );
  GTECH_XNOR4 U317 ( .A(n309), .B(n300), .C(n303), .D(n299), .Z(n335) );
  GTECH_XOR2 U318 ( .A(n321), .B(n336), .Z(n299) );
  GTECH_AND2 U319 ( .A(I_b[6]), .B(I_a[0]), .Z(n336) );
  GTECH_XOR3 U320 ( .A(n337), .B(n338), .C(n318), .Z(n321) );
  GTECH_NAND3 U321 ( .A(I_b[4]), .B(I_a[1]), .C(n339), .Z(n318) );
  GTECH_NOT U322 ( .A(n317), .Z(n338) );
  GTECH_NAND2 U323 ( .A(I_b[5]), .B(I_a[1]), .Z(n317) );
  GTECH_NOT U324 ( .A(n316), .Z(n337) );
  GTECH_NAND2 U325 ( .A(I_b[4]), .B(I_a[2]), .Z(n316) );
  GTECH_XOR3 U326 ( .A(n310), .B(n311), .C(n332), .Z(n303) );
  GTECH_OAI21 U327 ( .A(n340), .B(n341), .C(n342), .Z(n332) );
  GTECH_OAI21 U328 ( .A(n343), .B(n344), .C(n345), .Z(n342) );
  GTECH_NOT U329 ( .A(n346), .Z(n311) );
  GTECH_NAND2 U330 ( .A(I_a[5]), .B(I_b[1]), .Z(n346) );
  GTECH_NOT U331 ( .A(n330), .Z(n310) );
  GTECH_NAND2 U332 ( .A(I_a[6]), .B(I_b[0]), .Z(n330) );
  GTECH_ADD_ABC U333 ( .A(n347), .B(n348), .C(n349), .COUT(n300) );
  GTECH_NOT U334 ( .A(n350), .Z(n349) );
  GTECH_XOR3 U335 ( .A(n343), .B(n345), .C(n340), .Z(n348) );
  GTECH_NOT U336 ( .A(n344), .Z(n340) );
  GTECH_XOR3 U337 ( .A(n325), .B(n327), .C(n326), .Z(n309) );
  GTECH_OAI21 U338 ( .A(n351), .B(n352), .C(n353), .Z(n326) );
  GTECH_OAI21 U339 ( .A(n354), .B(n355), .C(n356), .Z(n353) );
  GTECH_NOT U340 ( .A(n355), .Z(n351) );
  GTECH_NOT U341 ( .A(n357), .Z(n327) );
  GTECH_NAND2 U342 ( .A(I_b[3]), .B(I_a[3]), .Z(n357) );
  GTECH_NOT U343 ( .A(n323), .Z(n325) );
  GTECH_NAND2 U344 ( .A(I_b[2]), .B(I_a[4]), .Z(n323) );
  GTECH_OA22 U345 ( .A(n306), .B(n307), .C(n358), .D(n305), .Z(n334) );
  GTECH_AND_NOT U346 ( .A(n306), .B(n359), .Z(n358) );
  GTECH_XOR3 U347 ( .A(n360), .B(n307), .C(n306), .Z(N145) );
  GTECH_XOR2 U348 ( .A(n361), .B(n339), .Z(n306) );
  GTECH_NOT U349 ( .A(n362), .Z(n339) );
  GTECH_NAND2 U350 ( .A(I_b[5]), .B(I_a[0]), .Z(n362) );
  GTECH_NAND2 U351 ( .A(I_b[4]), .B(I_a[1]), .Z(n361) );
  GTECH_NOT U352 ( .A(n359), .Z(n307) );
  GTECH_XOR2 U353 ( .A(n363), .B(n347), .Z(n359) );
  GTECH_ADD_ABC U354 ( .A(n364), .B(n365), .C(n366), .COUT(n347) );
  GTECH_XOR3 U355 ( .A(n367), .B(n368), .C(n369), .Z(n365) );
  GTECH_OA22 U356 ( .A(n370), .B(n371), .C(n372), .D(n373), .Z(n364) );
  GTECH_AND2 U357 ( .A(n372), .B(n373), .Z(n370) );
  GTECH_XNOR4 U358 ( .A(n345), .B(n344), .C(n350), .D(n343), .Z(n363) );
  GTECH_NOT U359 ( .A(n341), .Z(n343) );
  GTECH_NAND2 U360 ( .A(I_a[5]), .B(I_b[0]), .Z(n341) );
  GTECH_XOR3 U361 ( .A(n354), .B(n356), .C(n355), .Z(n350) );
  GTECH_OAI21 U362 ( .A(n374), .B(n375), .C(n376), .Z(n355) );
  GTECH_NOT U363 ( .A(n377), .Z(n356) );
  GTECH_NAND2 U364 ( .A(I_b[3]), .B(I_a[2]), .Z(n377) );
  GTECH_NOT U365 ( .A(n352), .Z(n354) );
  GTECH_NAND2 U366 ( .A(I_b[2]), .B(I_a[3]), .Z(n352) );
  GTECH_OAI21 U367 ( .A(n369), .B(n378), .C(n379), .Z(n344) );
  GTECH_OAI21 U368 ( .A(n367), .B(n380), .C(n368), .Z(n379) );
  GTECH_NOT U369 ( .A(n378), .Z(n367) );
  GTECH_NOT U370 ( .A(n380), .Z(n369) );
  GTECH_NOT U371 ( .A(n381), .Z(n345) );
  GTECH_NAND2 U372 ( .A(I_a[4]), .B(I_b[1]), .Z(n381) );
  GTECH_NOT U373 ( .A(n305), .Z(n360) );
  GTECH_NAND3 U374 ( .A(I_a[0]), .B(n382), .C(I_b[4]), .Z(n305) );
  GTECH_XOR2 U375 ( .A(n383), .B(n382), .Z(N144) );
  GTECH_XOR2 U376 ( .A(n384), .B(n385), .Z(n382) );
  GTECH_XNOR4 U377 ( .A(n368), .B(n380), .C(n378), .D(n366), .Z(n385) );
  GTECH_XOR3 U378 ( .A(n386), .B(n387), .C(n376), .Z(n366) );
  GTECH_NAND3 U379 ( .A(I_b[2]), .B(I_a[1]), .C(n388), .Z(n376) );
  GTECH_NOT U380 ( .A(n375), .Z(n387) );
  GTECH_NAND2 U381 ( .A(I_b[3]), .B(I_a[1]), .Z(n375) );
  GTECH_NOT U382 ( .A(n374), .Z(n386) );
  GTECH_NAND2 U383 ( .A(I_b[2]), .B(I_a[2]), .Z(n374) );
  GTECH_NAND2 U384 ( .A(I_a[4]), .B(I_b[0]), .Z(n378) );
  GTECH_OAI21 U385 ( .A(n389), .B(n390), .C(n391), .Z(n380) );
  GTECH_OAI21 U386 ( .A(n392), .B(n393), .C(n394), .Z(n391) );
  GTECH_NOT U387 ( .A(n393), .Z(n389) );
  GTECH_NOT U388 ( .A(n395), .Z(n368) );
  GTECH_NAND2 U389 ( .A(I_a[3]), .B(I_b[1]), .Z(n395) );
  GTECH_OA22 U390 ( .A(n372), .B(n373), .C(n396), .D(n371), .Z(n384) );
  GTECH_AND_NOT U391 ( .A(n372), .B(n397), .Z(n396) );
  GTECH_AND2 U392 ( .A(I_b[4]), .B(I_a[0]), .Z(n383) );
  GTECH_XOR3 U393 ( .A(n398), .B(n373), .C(n372), .Z(N143) );
  GTECH_XOR2 U394 ( .A(n399), .B(n388), .Z(n372) );
  GTECH_NOT U395 ( .A(n400), .Z(n388) );
  GTECH_NAND2 U396 ( .A(I_b[3]), .B(I_a[0]), .Z(n400) );
  GTECH_NAND2 U397 ( .A(I_b[2]), .B(I_a[1]), .Z(n399) );
  GTECH_NOT U398 ( .A(n397), .Z(n373) );
  GTECH_XOR3 U399 ( .A(n392), .B(n394), .C(n393), .Z(n397) );
  GTECH_OAI21 U400 ( .A(n401), .B(n402), .C(n403), .Z(n393) );
  GTECH_NOT U401 ( .A(n404), .Z(n394) );
  GTECH_NAND2 U402 ( .A(I_b[1]), .B(I_a[2]), .Z(n404) );
  GTECH_NOT U403 ( .A(n390), .Z(n392) );
  GTECH_NAND2 U404 ( .A(I_b[0]), .B(I_a[3]), .Z(n390) );
  GTECH_NOT U405 ( .A(n371), .Z(n398) );
  GTECH_NAND3 U406 ( .A(I_a[0]), .B(n405), .C(I_b[2]), .Z(n371) );
  GTECH_XOR2 U407 ( .A(n406), .B(n405), .Z(N142) );
  GTECH_NOT U408 ( .A(n407), .Z(n405) );
  GTECH_XOR3 U409 ( .A(n408), .B(n409), .C(n403), .Z(n407) );
  GTECH_NAND3 U410 ( .A(n410), .B(I_b[0]), .C(I_a[1]), .Z(n403) );
  GTECH_NOT U411 ( .A(n401), .Z(n409) );
  GTECH_NAND2 U412 ( .A(I_a[1]), .B(I_b[1]), .Z(n401) );
  GTECH_NOT U413 ( .A(n402), .Z(n408) );
  GTECH_NAND2 U414 ( .A(I_b[0]), .B(I_a[2]), .Z(n402) );
  GTECH_AND2 U415 ( .A(I_b[2]), .B(I_a[0]), .Z(n406) );
  GTECH_XOR2 U416 ( .A(n410), .B(n411), .Z(N141) );
  GTECH_AND2 U417 ( .A(I_a[1]), .B(I_b[0]), .Z(n411) );
  GTECH_NOT U418 ( .A(n412), .Z(n410) );
  GTECH_NAND2 U419 ( .A(I_a[0]), .B(I_b[1]), .Z(n412) );
  GTECH_AND2 U420 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

