
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n85) );
  GTECH_XNOR2 U78 ( .A(n84), .B(n90), .Z(N154) );
  GTECH_XNOR2 U79 ( .A(n91), .B(n92), .Z(n90) );
  GTECH_NOT U80 ( .A(n86), .Z(n92) );
  GTECH_XNOR2 U81 ( .A(n93), .B(n88), .Z(n86) );
  GTECH_NOT U82 ( .A(n94), .Z(n88) );
  GTECH_NAND2 U83 ( .A(I_b[7]), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U84 ( .A(n89), .Z(n93) );
  GTECH_OAI21 U85 ( .A(n95), .B(n96), .C(n97), .Z(n89) );
  GTECH_OAI21 U86 ( .A(n98), .B(n99), .C(n100), .Z(n97) );
  GTECH_NOT U87 ( .A(n87), .Z(n91) );
  GTECH_OAI2N2 U88 ( .A(n101), .B(n102), .C(n103), .D(n104), .Z(n87) );
  GTECH_NAND2 U89 ( .A(n101), .B(n102), .Z(n104) );
  GTECH_NOT U90 ( .A(n105), .Z(n84) );
  GTECH_NAND2 U91 ( .A(n106), .B(n107), .Z(n105) );
  GTECH_NOT U92 ( .A(n108), .Z(n106) );
  GTECH_XNOR2 U93 ( .A(n107), .B(n108), .Z(N153) );
  GTECH_XNOR3 U94 ( .A(n109), .B(n101), .C(n110), .Z(n108) );
  GTECH_NOT U95 ( .A(n103), .Z(n110) );
  GTECH_XNOR3 U96 ( .A(n98), .B(n100), .C(n95), .Z(n103) );
  GTECH_NOT U97 ( .A(n99), .Z(n95) );
  GTECH_OAI21 U98 ( .A(n111), .B(n112), .C(n113), .Z(n99) );
  GTECH_OAI21 U99 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_NOT U100 ( .A(n117), .Z(n100) );
  GTECH_NAND2 U101 ( .A(I_b[7]), .B(I_a[6]), .Z(n117) );
  GTECH_NOT U102 ( .A(n96), .Z(n98) );
  GTECH_NAND2 U103 ( .A(I_a[7]), .B(I_b[6]), .Z(n96) );
  GTECH_ADD_ABC U104 ( .A(n118), .B(n119), .C(n120), .COUT(n101) );
  GTECH_NOT U105 ( .A(n121), .Z(n120) );
  GTECH_XNOR2 U106 ( .A(n122), .B(n123), .Z(n119) );
  GTECH_NAND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n123) );
  GTECH_NOT U108 ( .A(n102), .Z(n109) );
  GTECH_NAND2 U109 ( .A(I_a[7]), .B(n124), .Z(n102) );
  GTECH_NOT U110 ( .A(n125), .Z(n107) );
  GTECH_NAND2 U111 ( .A(n126), .B(n127), .Z(n125) );
  GTECH_NOT U112 ( .A(n128), .Z(n127) );
  GTECH_XNOR2 U113 ( .A(n128), .B(n126), .Z(N152) );
  GTECH_XOR4 U114 ( .A(n122), .B(n129), .C(n121), .D(n118), .Z(n126) );
  GTECH_ADD_ABC U115 ( .A(n130), .B(n131), .C(n132), .COUT(n118) );
  GTECH_XNOR3 U116 ( .A(n133), .B(n134), .C(n135), .Z(n131) );
  GTECH_XNOR3 U117 ( .A(n114), .B(n116), .C(n111), .Z(n121) );
  GTECH_NOT U118 ( .A(n115), .Z(n111) );
  GTECH_OAI21 U119 ( .A(n136), .B(n137), .C(n138), .Z(n115) );
  GTECH_OAI21 U120 ( .A(n139), .B(n140), .C(n141), .Z(n138) );
  GTECH_NOT U121 ( .A(n142), .Z(n116) );
  GTECH_NAND2 U122 ( .A(I_b[7]), .B(I_a[5]), .Z(n142) );
  GTECH_NOT U123 ( .A(n112), .Z(n114) );
  GTECH_NAND2 U124 ( .A(I_b[6]), .B(I_a[6]), .Z(n112) );
  GTECH_AND2 U125 ( .A(I_a[7]), .B(I_b[5]), .Z(n129) );
  GTECH_NOT U126 ( .A(n124), .Z(n122) );
  GTECH_OAI21 U127 ( .A(n143), .B(n144), .C(n145), .Z(n124) );
  GTECH_OAI21 U128 ( .A(n133), .B(n135), .C(n134), .Z(n145) );
  GTECH_NOT U129 ( .A(n135), .Z(n143) );
  GTECH_ADD_ABC U130 ( .A(n146), .B(n147), .C(n148), .COUT(n128) );
  GTECH_OA22 U131 ( .A(n149), .B(n150), .C(n151), .D(n152), .Z(n147) );
  GTECH_OA21 U132 ( .A(n153), .B(n154), .C(n155), .Z(n146) );
  GTECH_XNOR3 U133 ( .A(n156), .B(n148), .C(n157), .Z(N151) );
  GTECH_OA21 U134 ( .A(n153), .B(n154), .C(n155), .Z(n157) );
  GTECH_OAI21 U135 ( .A(n158), .B(n159), .C(n160), .Z(n155) );
  GTECH_XOR4 U136 ( .A(n133), .B(n161), .C(n130), .D(n132), .Z(n148) );
  GTECH_NOT U137 ( .A(n162), .Z(n132) );
  GTECH_XNOR3 U138 ( .A(n139), .B(n141), .C(n136), .Z(n162) );
  GTECH_NOT U139 ( .A(n140), .Z(n136) );
  GTECH_OAI21 U140 ( .A(n163), .B(n164), .C(n165), .Z(n140) );
  GTECH_OAI21 U141 ( .A(n166), .B(n167), .C(n168), .Z(n165) );
  GTECH_NOT U142 ( .A(n169), .Z(n141) );
  GTECH_NAND2 U143 ( .A(I_b[7]), .B(I_a[4]), .Z(n169) );
  GTECH_NOT U144 ( .A(n137), .Z(n139) );
  GTECH_NAND2 U145 ( .A(I_b[6]), .B(I_a[5]), .Z(n137) );
  GTECH_ADD_ABC U146 ( .A(n170), .B(n171), .C(n172), .COUT(n130) );
  GTECH_NOT U147 ( .A(n173), .Z(n172) );
  GTECH_XNOR3 U148 ( .A(n174), .B(n175), .C(n176), .Z(n171) );
  GTECH_XNOR2 U149 ( .A(n134), .B(n135), .Z(n161) );
  GTECH_OAI21 U150 ( .A(n177), .B(n178), .C(n179), .Z(n135) );
  GTECH_OAI21 U151 ( .A(n174), .B(n176), .C(n175), .Z(n179) );
  GTECH_NOT U152 ( .A(n176), .Z(n177) );
  GTECH_NOT U153 ( .A(n180), .Z(n134) );
  GTECH_NAND2 U154 ( .A(I_a[6]), .B(I_b[5]), .Z(n180) );
  GTECH_NOT U155 ( .A(n144), .Z(n133) );
  GTECH_NAND2 U156 ( .A(I_a[7]), .B(I_b[4]), .Z(n144) );
  GTECH_OA22 U157 ( .A(n149), .B(n150), .C(n151), .D(n152), .Z(n156) );
  GTECH_NOT U158 ( .A(I_a[7]), .Z(n150) );
  GTECH_XNOR3 U159 ( .A(n153), .B(n158), .C(n160), .Z(N150) );
  GTECH_XOR4 U160 ( .A(n174), .B(n181), .C(n173), .D(n170), .Z(n160) );
  GTECH_ADD_ABC U161 ( .A(n182), .B(n183), .C(n184), .COUT(n170) );
  GTECH_NOT U162 ( .A(n185), .Z(n184) );
  GTECH_XNOR3 U163 ( .A(n186), .B(n187), .C(n188), .Z(n183) );
  GTECH_XNOR3 U164 ( .A(n166), .B(n168), .C(n163), .Z(n173) );
  GTECH_NOT U165 ( .A(n167), .Z(n163) );
  GTECH_OAI21 U166 ( .A(n189), .B(n190), .C(n191), .Z(n167) );
  GTECH_OAI21 U167 ( .A(n192), .B(n193), .C(n194), .Z(n191) );
  GTECH_NOT U168 ( .A(n195), .Z(n168) );
  GTECH_NAND2 U169 ( .A(I_b[7]), .B(I_a[3]), .Z(n195) );
  GTECH_NOT U170 ( .A(n164), .Z(n166) );
  GTECH_NAND2 U171 ( .A(I_b[6]), .B(I_a[4]), .Z(n164) );
  GTECH_XNOR2 U172 ( .A(n175), .B(n176), .Z(n181) );
  GTECH_OAI21 U173 ( .A(n196), .B(n197), .C(n198), .Z(n176) );
  GTECH_OAI21 U174 ( .A(n186), .B(n188), .C(n187), .Z(n198) );
  GTECH_NOT U175 ( .A(n188), .Z(n196) );
  GTECH_NOT U176 ( .A(n199), .Z(n175) );
  GTECH_NAND2 U177 ( .A(I_a[5]), .B(I_b[5]), .Z(n199) );
  GTECH_NOT U178 ( .A(n178), .Z(n174) );
  GTECH_NAND2 U179 ( .A(I_a[6]), .B(I_b[4]), .Z(n178) );
  GTECH_NOT U180 ( .A(n154), .Z(n158) );
  GTECH_XNOR2 U181 ( .A(n151), .B(n152), .Z(n154) );
  GTECH_XNOR2 U182 ( .A(n149), .B(n200), .Z(n152) );
  GTECH_NAND2 U183 ( .A(I_a[7]), .B(I_b[3]), .Z(n200) );
  GTECH_OA21 U184 ( .A(n201), .B(n202), .C(n203), .Z(n149) );
  GTECH_OAI21 U185 ( .A(n204), .B(n205), .C(n206), .Z(n203) );
  GTECH_AOI2N2 U186 ( .A(n207), .B(n208), .C(n209), .D(n210), .Z(n151) );
  GTECH_NAND2 U187 ( .A(n209), .B(n210), .Z(n208) );
  GTECH_NOT U188 ( .A(n159), .Z(n153) );
  GTECH_OAI2N2 U189 ( .A(n211), .B(n212), .C(n213), .D(n214), .Z(n159) );
  GTECH_NAND2 U190 ( .A(n211), .B(n212), .Z(n214) );
  GTECH_XNOR3 U191 ( .A(n211), .B(n215), .C(n213), .Z(N149) );
  GTECH_XOR4 U192 ( .A(n186), .B(n216), .C(n185), .D(n182), .Z(n213) );
  GTECH_ADD_ABC U193 ( .A(n217), .B(n218), .C(n219), .COUT(n182) );
  GTECH_XNOR3 U194 ( .A(n220), .B(n221), .C(n222), .Z(n218) );
  GTECH_OA21 U195 ( .A(n223), .B(n224), .C(n225), .Z(n217) );
  GTECH_XNOR3 U196 ( .A(n192), .B(n194), .C(n189), .Z(n185) );
  GTECH_NOT U197 ( .A(n193), .Z(n189) );
  GTECH_OAI21 U198 ( .A(n226), .B(n227), .C(n228), .Z(n193) );
  GTECH_NOT U199 ( .A(n229), .Z(n194) );
  GTECH_NAND2 U200 ( .A(I_b[7]), .B(I_a[2]), .Z(n229) );
  GTECH_NOT U201 ( .A(n190), .Z(n192) );
  GTECH_NAND2 U202 ( .A(I_b[6]), .B(I_a[3]), .Z(n190) );
  GTECH_XNOR2 U203 ( .A(n187), .B(n188), .Z(n216) );
  GTECH_OAI21 U204 ( .A(n230), .B(n231), .C(n232), .Z(n188) );
  GTECH_OAI21 U205 ( .A(n220), .B(n222), .C(n221), .Z(n232) );
  GTECH_NOT U206 ( .A(n222), .Z(n230) );
  GTECH_NOT U207 ( .A(n233), .Z(n187) );
  GTECH_NAND2 U208 ( .A(I_b[5]), .B(I_a[4]), .Z(n233) );
  GTECH_NOT U209 ( .A(n197), .Z(n186) );
  GTECH_NAND2 U210 ( .A(I_a[5]), .B(I_b[4]), .Z(n197) );
  GTECH_NOT U211 ( .A(n212), .Z(n215) );
  GTECH_XNOR3 U212 ( .A(n234), .B(n209), .C(n235), .Z(n212) );
  GTECH_NOT U213 ( .A(n207), .Z(n235) );
  GTECH_XNOR3 U214 ( .A(n204), .B(n206), .C(n201), .Z(n207) );
  GTECH_NOT U215 ( .A(n205), .Z(n201) );
  GTECH_OAI21 U216 ( .A(n236), .B(n237), .C(n238), .Z(n205) );
  GTECH_OAI21 U217 ( .A(n239), .B(n240), .C(n241), .Z(n238) );
  GTECH_NOT U218 ( .A(n242), .Z(n206) );
  GTECH_NAND2 U219 ( .A(I_a[6]), .B(I_b[3]), .Z(n242) );
  GTECH_NOT U220 ( .A(n202), .Z(n204) );
  GTECH_NAND2 U221 ( .A(I_a[7]), .B(I_b[2]), .Z(n202) );
  GTECH_ADD_ABC U222 ( .A(n243), .B(n244), .C(n245), .COUT(n209) );
  GTECH_XNOR2 U223 ( .A(n246), .B(n247), .Z(n244) );
  GTECH_NAND2 U224 ( .A(I_a[7]), .B(I_b[1]), .Z(n247) );
  GTECH_NOT U225 ( .A(n210), .Z(n234) );
  GTECH_NAND2 U226 ( .A(I_a[7]), .B(n248), .Z(n210) );
  GTECH_ADD_ABC U227 ( .A(n249), .B(n250), .C(n251), .COUT(n211) );
  GTECH_XNOR3 U228 ( .A(n243), .B(n252), .C(n253), .Z(n250) );
  GTECH_XOR4 U229 ( .A(n243), .B(n251), .C(n254), .D(n249), .Z(N148) );
  GTECH_ADD_ABC U230 ( .A(n255), .B(n256), .C(n257), .COUT(n249) );
  GTECH_NOT U231 ( .A(n258), .Z(n257) );
  GTECH_XNOR3 U232 ( .A(n259), .B(n260), .C(n261), .Z(n256) );
  GTECH_XNOR2 U233 ( .A(n252), .B(n245), .Z(n254) );
  GTECH_NOT U234 ( .A(n253), .Z(n245) );
  GTECH_XNOR3 U235 ( .A(n239), .B(n241), .C(n236), .Z(n253) );
  GTECH_NOT U236 ( .A(n240), .Z(n236) );
  GTECH_OAI21 U237 ( .A(n262), .B(n263), .C(n264), .Z(n240) );
  GTECH_OAI21 U238 ( .A(n265), .B(n266), .C(n267), .Z(n264) );
  GTECH_NOT U239 ( .A(n268), .Z(n241) );
  GTECH_NAND2 U240 ( .A(I_a[5]), .B(I_b[3]), .Z(n268) );
  GTECH_NOT U241 ( .A(n237), .Z(n239) );
  GTECH_NAND2 U242 ( .A(I_a[6]), .B(I_b[2]), .Z(n237) );
  GTECH_XNOR2 U243 ( .A(n246), .B(n269), .Z(n252) );
  GTECH_NAND2 U244 ( .A(I_a[7]), .B(I_b[1]), .Z(n269) );
  GTECH_NOT U245 ( .A(n248), .Z(n246) );
  GTECH_OAI21 U246 ( .A(n270), .B(n271), .C(n272), .Z(n248) );
  GTECH_OAI21 U247 ( .A(n273), .B(n274), .C(n275), .Z(n272) );
  GTECH_XOR4 U248 ( .A(n220), .B(n276), .C(n277), .D(n219), .Z(n251) );
  GTECH_XNOR3 U249 ( .A(n278), .B(n279), .C(n280), .Z(n219) );
  GTECH_NOT U250 ( .A(n228), .Z(n280) );
  GTECH_NAND3 U251 ( .A(I_b[6]), .B(I_a[1]), .C(n281), .Z(n228) );
  GTECH_NOT U252 ( .A(n227), .Z(n279) );
  GTECH_NAND2 U253 ( .A(I_b[7]), .B(I_a[1]), .Z(n227) );
  GTECH_NOT U254 ( .A(n226), .Z(n278) );
  GTECH_NAND2 U255 ( .A(I_b[6]), .B(I_a[2]), .Z(n226) );
  GTECH_OA21 U256 ( .A(n223), .B(n224), .C(n225), .Z(n277) );
  GTECH_OAI21 U257 ( .A(n282), .B(n283), .C(n284), .Z(n225) );
  GTECH_XNOR2 U258 ( .A(n221), .B(n222), .Z(n276) );
  GTECH_OAI21 U259 ( .A(n285), .B(n286), .C(n287), .Z(n222) );
  GTECH_OAI21 U260 ( .A(n288), .B(n289), .C(n290), .Z(n287) );
  GTECH_NOT U261 ( .A(n291), .Z(n221) );
  GTECH_NAND2 U262 ( .A(I_b[5]), .B(I_a[3]), .Z(n291) );
  GTECH_NOT U263 ( .A(n231), .Z(n220) );
  GTECH_NAND2 U264 ( .A(I_b[4]), .B(I_a[4]), .Z(n231) );
  GTECH_ADD_ABC U265 ( .A(n259), .B(n292), .C(n293), .COUT(n243) );
  GTECH_NOT U266 ( .A(n261), .Z(n293) );
  GTECH_XNOR3 U267 ( .A(n273), .B(n275), .C(n274), .Z(n292) );
  GTECH_XOR4 U268 ( .A(n259), .B(n294), .C(n258), .D(n255), .Z(N147) );
  GTECH_ADD_ABC U269 ( .A(n295), .B(n296), .C(n297), .COUT(n255) );
  GTECH_XNOR3 U270 ( .A(n298), .B(n299), .C(n300), .Z(n296) );
  GTECH_OA21 U271 ( .A(n301), .B(n302), .C(n303), .Z(n295) );
  GTECH_XNOR3 U272 ( .A(n284), .B(n224), .C(n283), .Z(n258) );
  GTECH_NOT U273 ( .A(n223), .Z(n283) );
  GTECH_XNOR2 U274 ( .A(n281), .B(n304), .Z(n223) );
  GTECH_AND2 U275 ( .A(I_b[6]), .B(I_a[1]), .Z(n304) );
  GTECH_NOT U276 ( .A(n305), .Z(n281) );
  GTECH_NAND2 U277 ( .A(I_b[7]), .B(I_a[0]), .Z(n305) );
  GTECH_NOT U278 ( .A(n282), .Z(n224) );
  GTECH_XNOR3 U279 ( .A(n288), .B(n290), .C(n285), .Z(n282) );
  GTECH_NOT U280 ( .A(n289), .Z(n285) );
  GTECH_OAI21 U281 ( .A(n306), .B(n307), .C(n308), .Z(n289) );
  GTECH_NOT U282 ( .A(n309), .Z(n290) );
  GTECH_NAND2 U283 ( .A(I_b[5]), .B(I_a[2]), .Z(n309) );
  GTECH_NOT U284 ( .A(n286), .Z(n288) );
  GTECH_NAND2 U285 ( .A(I_b[4]), .B(I_a[3]), .Z(n286) );
  GTECH_NOT U286 ( .A(n310), .Z(n284) );
  GTECH_NAND3 U287 ( .A(I_a[0]), .B(n311), .C(I_b[6]), .Z(n310) );
  GTECH_XNOR2 U288 ( .A(n260), .B(n261), .Z(n294) );
  GTECH_XNOR3 U289 ( .A(n265), .B(n267), .C(n262), .Z(n261) );
  GTECH_NOT U290 ( .A(n266), .Z(n262) );
  GTECH_OAI21 U291 ( .A(n312), .B(n313), .C(n314), .Z(n266) );
  GTECH_OAI21 U292 ( .A(n315), .B(n316), .C(n317), .Z(n314) );
  GTECH_NOT U293 ( .A(n318), .Z(n267) );
  GTECH_NAND2 U294 ( .A(I_b[3]), .B(I_a[4]), .Z(n318) );
  GTECH_NOT U295 ( .A(n263), .Z(n265) );
  GTECH_NAND2 U296 ( .A(I_a[5]), .B(I_b[2]), .Z(n263) );
  GTECH_NOT U297 ( .A(n319), .Z(n260) );
  GTECH_XNOR3 U298 ( .A(n273), .B(n275), .C(n270), .Z(n319) );
  GTECH_NOT U299 ( .A(n274), .Z(n270) );
  GTECH_OAI21 U300 ( .A(n320), .B(n321), .C(n322), .Z(n274) );
  GTECH_OAI21 U301 ( .A(n323), .B(n324), .C(n325), .Z(n322) );
  GTECH_NOT U302 ( .A(n326), .Z(n275) );
  GTECH_NAND2 U303 ( .A(I_a[6]), .B(I_b[1]), .Z(n326) );
  GTECH_NOT U304 ( .A(n271), .Z(n273) );
  GTECH_NAND2 U305 ( .A(I_a[7]), .B(I_b[0]), .Z(n271) );
  GTECH_ADD_ABC U306 ( .A(n298), .B(n327), .C(n328), .COUT(n259) );
  GTECH_NOT U307 ( .A(n300), .Z(n328) );
  GTECH_XNOR3 U308 ( .A(n323), .B(n325), .C(n324), .Z(n327) );
  GTECH_XOR4 U309 ( .A(n298), .B(n329), .C(n330), .D(n297), .Z(N146) );
  GTECH_XNOR2 U310 ( .A(n331), .B(n311), .Z(n297) );
  GTECH_NOT U311 ( .A(n332), .Z(n311) );
  GTECH_XNOR3 U312 ( .A(n333), .B(n334), .C(n335), .Z(n332) );
  GTECH_NOT U313 ( .A(n308), .Z(n335) );
  GTECH_NAND3 U314 ( .A(I_b[4]), .B(I_a[1]), .C(n336), .Z(n308) );
  GTECH_NOT U315 ( .A(n307), .Z(n334) );
  GTECH_NAND2 U316 ( .A(I_b[5]), .B(I_a[1]), .Z(n307) );
  GTECH_NOT U317 ( .A(n306), .Z(n333) );
  GTECH_NAND2 U318 ( .A(I_b[4]), .B(I_a[2]), .Z(n306) );
  GTECH_AND2 U319 ( .A(I_b[6]), .B(I_a[0]), .Z(n331) );
  GTECH_OAI21 U320 ( .A(n301), .B(n302), .C(n303), .Z(n330) );
  GTECH_OAI21 U321 ( .A(n337), .B(n338), .C(n339), .Z(n303) );
  GTECH_XNOR2 U322 ( .A(n299), .B(n300), .Z(n329) );
  GTECH_XNOR3 U323 ( .A(n315), .B(n317), .C(n312), .Z(n300) );
  GTECH_NOT U324 ( .A(n316), .Z(n312) );
  GTECH_OAI21 U325 ( .A(n340), .B(n341), .C(n342), .Z(n316) );
  GTECH_OAI21 U326 ( .A(n343), .B(n344), .C(n345), .Z(n342) );
  GTECH_NOT U327 ( .A(n346), .Z(n317) );
  GTECH_NAND2 U328 ( .A(I_b[3]), .B(I_a[3]), .Z(n346) );
  GTECH_NOT U329 ( .A(n313), .Z(n315) );
  GTECH_NAND2 U330 ( .A(I_b[2]), .B(I_a[4]), .Z(n313) );
  GTECH_NOT U331 ( .A(n347), .Z(n299) );
  GTECH_XNOR3 U332 ( .A(n323), .B(n325), .C(n320), .Z(n347) );
  GTECH_NOT U333 ( .A(n324), .Z(n320) );
  GTECH_OAI21 U334 ( .A(n348), .B(n349), .C(n350), .Z(n324) );
  GTECH_OAI21 U335 ( .A(n351), .B(n352), .C(n353), .Z(n350) );
  GTECH_NOT U336 ( .A(n352), .Z(n348) );
  GTECH_NOT U337 ( .A(n354), .Z(n325) );
  GTECH_NAND2 U338 ( .A(I_a[5]), .B(I_b[1]), .Z(n354) );
  GTECH_NOT U339 ( .A(n321), .Z(n323) );
  GTECH_NAND2 U340 ( .A(I_a[6]), .B(I_b[0]), .Z(n321) );
  GTECH_ADD_ABC U341 ( .A(n355), .B(n356), .C(n357), .COUT(n298) );
  GTECH_NOT U342 ( .A(n358), .Z(n357) );
  GTECH_XNOR3 U343 ( .A(n351), .B(n353), .C(n352), .Z(n356) );
  GTECH_XNOR3 U344 ( .A(n339), .B(n302), .C(n338), .Z(N145) );
  GTECH_NOT U345 ( .A(n301), .Z(n338) );
  GTECH_XNOR2 U346 ( .A(n336), .B(n359), .Z(n301) );
  GTECH_AND2 U347 ( .A(I_b[4]), .B(I_a[1]), .Z(n359) );
  GTECH_NOT U348 ( .A(n360), .Z(n336) );
  GTECH_NAND2 U349 ( .A(I_b[5]), .B(I_a[0]), .Z(n360) );
  GTECH_NOT U350 ( .A(n337), .Z(n302) );
  GTECH_XOR4 U351 ( .A(n351), .B(n361), .C(n358), .D(n355), .Z(n337) );
  GTECH_ADD_ABC U352 ( .A(n362), .B(n363), .C(n364), .COUT(n355) );
  GTECH_XNOR3 U353 ( .A(n365), .B(n366), .C(n367), .Z(n363) );
  GTECH_OA21 U354 ( .A(n368), .B(n369), .C(n370), .Z(n362) );
  GTECH_XNOR3 U355 ( .A(n343), .B(n345), .C(n340), .Z(n358) );
  GTECH_NOT U356 ( .A(n344), .Z(n340) );
  GTECH_OAI21 U357 ( .A(n371), .B(n372), .C(n373), .Z(n344) );
  GTECH_NOT U358 ( .A(n374), .Z(n345) );
  GTECH_NAND2 U359 ( .A(I_b[3]), .B(I_a[2]), .Z(n374) );
  GTECH_NOT U360 ( .A(n341), .Z(n343) );
  GTECH_NAND2 U361 ( .A(I_b[2]), .B(I_a[3]), .Z(n341) );
  GTECH_XNOR2 U362 ( .A(n353), .B(n352), .Z(n361) );
  GTECH_OAI21 U363 ( .A(n375), .B(n376), .C(n377), .Z(n352) );
  GTECH_OAI21 U364 ( .A(n365), .B(n367), .C(n366), .Z(n377) );
  GTECH_NOT U365 ( .A(n367), .Z(n375) );
  GTECH_NOT U366 ( .A(n378), .Z(n353) );
  GTECH_NAND2 U367 ( .A(I_a[4]), .B(I_b[1]), .Z(n378) );
  GTECH_NOT U368 ( .A(n349), .Z(n351) );
  GTECH_NAND2 U369 ( .A(I_a[5]), .B(I_b[0]), .Z(n349) );
  GTECH_NOT U370 ( .A(n379), .Z(n339) );
  GTECH_NAND3 U371 ( .A(I_a[0]), .B(n380), .C(I_b[4]), .Z(n379) );
  GTECH_NOT U372 ( .A(n381), .Z(n380) );
  GTECH_XNOR2 U373 ( .A(n382), .B(n381), .Z(N144) );
  GTECH_XOR4 U374 ( .A(n365), .B(n383), .C(n384), .D(n364), .Z(n381) );
  GTECH_XNOR3 U375 ( .A(n385), .B(n386), .C(n387), .Z(n364) );
  GTECH_NOT U376 ( .A(n373), .Z(n387) );
  GTECH_NAND3 U377 ( .A(I_b[2]), .B(I_a[1]), .C(n388), .Z(n373) );
  GTECH_NOT U378 ( .A(n372), .Z(n386) );
  GTECH_NAND2 U379 ( .A(I_b[3]), .B(I_a[1]), .Z(n372) );
  GTECH_NOT U380 ( .A(n371), .Z(n385) );
  GTECH_NAND2 U381 ( .A(I_b[2]), .B(I_a[2]), .Z(n371) );
  GTECH_OA21 U382 ( .A(n368), .B(n369), .C(n370), .Z(n384) );
  GTECH_OAI21 U383 ( .A(n389), .B(n390), .C(n391), .Z(n370) );
  GTECH_XNOR2 U384 ( .A(n366), .B(n367), .Z(n383) );
  GTECH_OAI21 U385 ( .A(n392), .B(n393), .C(n394), .Z(n367) );
  GTECH_OAI21 U386 ( .A(n395), .B(n396), .C(n397), .Z(n394) );
  GTECH_NOT U387 ( .A(n398), .Z(n366) );
  GTECH_NAND2 U388 ( .A(I_a[3]), .B(I_b[1]), .Z(n398) );
  GTECH_NOT U389 ( .A(n376), .Z(n365) );
  GTECH_NAND2 U390 ( .A(I_a[4]), .B(I_b[0]), .Z(n376) );
  GTECH_AND2 U391 ( .A(I_b[4]), .B(I_a[0]), .Z(n382) );
  GTECH_XNOR3 U392 ( .A(n391), .B(n369), .C(n390), .Z(N143) );
  GTECH_NOT U393 ( .A(n368), .Z(n390) );
  GTECH_XNOR2 U394 ( .A(n388), .B(n399), .Z(n368) );
  GTECH_AND2 U395 ( .A(I_b[2]), .B(I_a[1]), .Z(n399) );
  GTECH_NOT U396 ( .A(n400), .Z(n388) );
  GTECH_NAND2 U397 ( .A(I_b[3]), .B(I_a[0]), .Z(n400) );
  GTECH_NOT U398 ( .A(n389), .Z(n369) );
  GTECH_XNOR3 U399 ( .A(n395), .B(n397), .C(n392), .Z(n389) );
  GTECH_NOT U400 ( .A(n396), .Z(n392) );
  GTECH_OAI21 U401 ( .A(n401), .B(n402), .C(n403), .Z(n396) );
  GTECH_NOT U402 ( .A(n404), .Z(n397) );
  GTECH_NAND2 U403 ( .A(I_b[1]), .B(I_a[2]), .Z(n404) );
  GTECH_NOT U404 ( .A(n393), .Z(n395) );
  GTECH_NAND2 U405 ( .A(I_b[0]), .B(I_a[3]), .Z(n393) );
  GTECH_NOT U406 ( .A(n405), .Z(n391) );
  GTECH_NAND3 U407 ( .A(I_a[0]), .B(n406), .C(I_b[2]), .Z(n405) );
  GTECH_NOT U408 ( .A(n407), .Z(n406) );
  GTECH_XNOR2 U409 ( .A(n408), .B(n407), .Z(N142) );
  GTECH_XNOR3 U410 ( .A(n409), .B(n410), .C(n411), .Z(n407) );
  GTECH_NOT U411 ( .A(n403), .Z(n411) );
  GTECH_NAND3 U412 ( .A(n412), .B(I_b[0]), .C(I_a[1]), .Z(n403) );
  GTECH_NOT U413 ( .A(n401), .Z(n410) );
  GTECH_NAND2 U414 ( .A(I_a[1]), .B(I_b[1]), .Z(n401) );
  GTECH_NOT U415 ( .A(n402), .Z(n409) );
  GTECH_NAND2 U416 ( .A(I_b[0]), .B(I_a[2]), .Z(n402) );
  GTECH_AND2 U417 ( .A(I_b[2]), .B(I_a[0]), .Z(n408) );
  GTECH_XNOR2 U418 ( .A(n412), .B(n413), .Z(N141) );
  GTECH_NAND2 U419 ( .A(I_a[1]), .B(I_b[0]), .Z(n413) );
  GTECH_NOT U420 ( .A(n414), .Z(n412) );
  GTECH_NAND2 U421 ( .A(I_a[0]), .B(I_b[1]), .Z(n414) );
  GTECH_AND2 U422 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

