
module shift_add_multiplier ( clk, rst, D, Q, out );
  input [7:0] D;
  input [7:0] Q;
  output [15:0] out;
  input clk, rst;
  wire   load_cmd, add_cmd, shift_cmd, out_cmd, lsb, shifter_N24, shifter_N23,
         shifter_N22, shifter_N21, shifter_N20, shifter_N19, shifter_N18,
         shifter_N17, shifter_N16, shifter_N15, shifter_N14, shifter_N13,
         shifter_N12, shifter_N11, shifter_N10, shifter_N9, shifter_N8,
         shifter_N7, shifter_N6, shifter_add_temp, shifter_temp_1_,
         shifter_temp_2_, shifter_temp_3_, shifter_temp_4_, shifter_temp_5_,
         shifter_temp_6_, shifter_temp_7_, controller_N102, controller_N98,
         controller_N97, controller_N96, controller_N95, controller_N94,
         controller_N93, controller_N92, controller_N91, controller_N90,
         controller_N83, controller_N82, controller_N81, controller_N80,
         controller_N79, controller_N78, controller_N77, controller_N76,
         controller_N75, controller_N74, controller_N73, controller_N72,
         controller_N71, controller_N70, controller_N69, controller_N68,
         controller_N67, controller_N66, controller_N65, controller_N64,
         controller_N63, controller_N62, controller_N61, controller_N60,
         controller_N59, controller_N58, controller_N57, controller_N56,
         controller_N55, controller_N54, controller_N53, controller_N52,
         controller_count_0_, controller_count_1_, controller_count_2_,
         controller_count_3_, controller_count_4_, controller_count_5_,
         controller_count_6_, controller_count_7_, controller_count_8_,
         controller_count_9_, controller_count_10_, controller_count_11_,
         controller_count_12_, controller_count_13_, controller_count_14_,
         controller_count_15_, controller_count_16_, controller_count_17_,
         controller_count_18_, controller_count_19_, controller_count_20_,
         controller_count_21_, controller_count_22_, controller_count_23_,
         controller_count_24_, controller_count_25_, controller_count_26_,
         controller_count_27_, controller_count_28_, controller_count_29_,
         controller_count_30_, controller_count_31_, controller_state_0_,
         controller_state_1_, controller_state_2_, controller_start, n8, n11,
         n12, n13, n14, n15, n16, n17, n18, n127, n129, n132, n43, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370;
  wire   [7:0] A;

  GTECH_FJK2S controller_count_reg_31_ ( .J(n43), .K(n43), .TI(controller_N83), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_31_), 
        .QN(n153) );
  GTECH_FJK2S controller_count_reg_30_ ( .J(n43), .K(n43), .TI(controller_N82), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_30_), 
        .QN(n152) );
  GTECH_FJK3 controller_start_reg ( .J(n43), .K(controller_N97), .CP(clk), 
        .CD(n127), .SD(n132), .Q(controller_start), .QN(n129) );
  GTECH_FJK2S controller_state_reg_0_ ( .J(n43), .K(n43), .TI(controller_N93), 
        .TE(controller_N95), .CP(clk), .CD(n132), .Q(controller_state_0_), 
        .QN(n138) );
  GTECH_FJK2S controller_state_reg_1_ ( .J(n43), .K(n43), .TI(controller_N94), 
        .TE(controller_N95), .CP(clk), .CD(n132), .Q(controller_state_1_), 
        .QN(n8) );
  GTECH_FJK2S controller_state_reg_2_ ( .J(n43), .K(n43), .TI(controller_N96), 
        .TE(controller_N95), .CP(clk), .CD(n132), .Q(controller_state_2_), 
        .QN(n139) );
  GTECH_FJK2S controller_count_reg_29_ ( .J(n43), .K(n43), .TI(controller_N81), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_29_), 
        .QN(n151) );
  GTECH_FJK2S controller_count_reg_28_ ( .J(n43), .K(n43), .TI(controller_N80), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_28_), 
        .QN(n150) );
  GTECH_FJK2S controller_count_reg_27_ ( .J(n43), .K(n43), .TI(controller_N79), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_27_), 
        .QN(n149) );
  GTECH_FJK2S controller_count_reg_26_ ( .J(n43), .K(n43), .TI(controller_N78), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_26_), 
        .QN(n148) );
  GTECH_FJK2S controller_count_reg_25_ ( .J(n43), .K(n43), .TI(controller_N77), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_25_), 
        .QN(n147) );
  GTECH_FJK2S controller_count_reg_24_ ( .J(n43), .K(n43), .TI(controller_N76), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_24_), 
        .QN(n146) );
  GTECH_FJK2S controller_count_reg_23_ ( .J(n43), .K(n43), .TI(controller_N75), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_23_), 
        .QN(n145) );
  GTECH_FJK2S controller_count_reg_22_ ( .J(n43), .K(n43), .TI(controller_N74), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_22_), 
        .QN(n144) );
  GTECH_FJK2S controller_count_reg_21_ ( .J(n43), .K(n43), .TI(controller_N73), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_21_), 
        .QN(n143) );
  GTECH_FJK2S controller_count_reg_20_ ( .J(n43), .K(n43), .TI(controller_N72), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_20_), 
        .QN(n142) );
  GTECH_FJK2S controller_count_reg_19_ ( .J(n43), .K(n43), .TI(controller_N71), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_19_), 
        .QN(n141) );
  GTECH_FJK2S controller_count_reg_18_ ( .J(n43), .K(n43), .TI(controller_N70), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_18_), 
        .QN(n140) );
  GTECH_FJK2S controller_count_reg_17_ ( .J(n43), .K(n43), .TI(controller_N69), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_17_), 
        .QN(n171) );
  GTECH_FJK2S controller_count_reg_16_ ( .J(n43), .K(n43), .TI(controller_N68), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_16_), 
        .QN(n170) );
  GTECH_FJK2S controller_count_reg_15_ ( .J(n43), .K(n43), .TI(controller_N67), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_15_), 
        .QN(n169) );
  GTECH_FJK2S controller_count_reg_14_ ( .J(n43), .K(n43), .TI(controller_N66), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_14_), 
        .QN(n168) );
  GTECH_FJK2S controller_count_reg_13_ ( .J(n43), .K(n43), .TI(controller_N65), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_13_), 
        .QN(n167) );
  GTECH_FJK2S controller_count_reg_12_ ( .J(n43), .K(n43), .TI(controller_N64), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_12_), 
        .QN(n166) );
  GTECH_FJK2S controller_count_reg_11_ ( .J(n43), .K(n43), .TI(controller_N63), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_11_), 
        .QN(n165) );
  GTECH_FJK2S controller_count_reg_10_ ( .J(n43), .K(n43), .TI(controller_N62), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_10_), 
        .QN(n164) );
  GTECH_FJK2S controller_count_reg_9_ ( .J(n43), .K(n43), .TI(controller_N61), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_9_), 
        .QN(n163) );
  GTECH_FJK2S controller_count_reg_8_ ( .J(n43), .K(n43), .TI(controller_N60), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_8_), 
        .QN(n162) );
  GTECH_FJK2S controller_count_reg_7_ ( .J(n43), .K(n43), .TI(controller_N59), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_7_), 
        .QN(n161) );
  GTECH_FJK2S controller_count_reg_6_ ( .J(n43), .K(n43), .TI(controller_N58), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_6_), 
        .QN(n160) );
  GTECH_FJK2S controller_count_reg_5_ ( .J(n43), .K(n43), .TI(controller_N57), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_5_), 
        .QN(n159) );
  GTECH_FJK2S controller_count_reg_4_ ( .J(n43), .K(n43), .TI(controller_N56), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_4_), 
        .QN(n158) );
  GTECH_FJK2S controller_count_reg_3_ ( .J(n43), .K(n43), .TI(controller_N55), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_3_), 
        .QN(n157) );
  GTECH_FJK2S controller_count_reg_2_ ( .J(n43), .K(n43), .TI(controller_N54), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_2_), 
        .QN(n156) );
  GTECH_FJK2S controller_count_reg_1_ ( .J(n43), .K(n43), .TI(controller_N53), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_1_), 
        .QN(n155) );
  GTECH_FJK2S controller_count_reg_0_ ( .J(n43), .K(n43), .TI(controller_N52), 
        .TE(controller_N98), .CP(clk), .CD(n132), .Q(controller_count_0_), 
        .QN(n154) );
  GTECH_FJK1S controller_shift_cmd_reg ( .J(n43), .K(n43), .TI(controller_N98), 
        .TE(controller_N102), .CP(clk), .Q(shift_cmd) );
  GTECH_FJK1S controller_add_cmd_reg ( .J(n43), .K(n43), .TI(controller_N91), 
        .TE(controller_N102), .CP(clk), .Q(add_cmd), .QN(n135) );
  GTECH_FJK1S controller_load_cmd_reg ( .J(n43), .K(n43), .TI(controller_N90), 
        .TE(controller_N102), .CP(clk), .Q(load_cmd), .QN(n136) );
  GTECH_FJK2S shifter_add_temp_reg ( .J(n43), .K(n43), .TI(shifter_N24), .TE(
        shifter_N23), .CP(clk), .CD(n132), .Q(shifter_add_temp) );
  GTECH_FJK2S shifter_temp_reg_8_ ( .J(n43), .K(n43), .TI(shifter_N14), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(A[0]), .QN(n11) );
  GTECH_FJK2S shifter_temp_reg_15_ ( .J(n43), .K(n43), .TI(shifter_N21), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(A[7]), .QN(n12) );
  GTECH_FJK2S shifter_temp_reg_14_ ( .J(n43), .K(n43), .TI(shifter_N20), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(A[6]), .QN(n13) );
  GTECH_FJK2S shifter_temp_reg_13_ ( .J(n43), .K(n43), .TI(shifter_N19), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(A[5]), .QN(n14) );
  GTECH_FJK2S shifter_temp_reg_12_ ( .J(n43), .K(n43), .TI(shifter_N18), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(A[4]), .QN(n15) );
  GTECH_FJK2S shifter_temp_reg_11_ ( .J(n43), .K(n43), .TI(shifter_N17), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(A[3]), .QN(n16) );
  GTECH_FJK2S shifter_temp_reg_10_ ( .J(n43), .K(n43), .TI(shifter_N16), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(A[2]), .QN(n17) );
  GTECH_FJK2S shifter_temp_reg_9_ ( .J(n43), .K(n43), .TI(shifter_N15), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(A[1]), .QN(n18) );
  GTECH_FJK2S shifter_temp_reg_7_ ( .J(n43), .K(n43), .TI(shifter_N13), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(shifter_temp_7_) );
  GTECH_FJK2S shifter_temp_reg_6_ ( .J(n43), .K(n43), .TI(shifter_N12), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(shifter_temp_6_) );
  GTECH_FJK2S shifter_temp_reg_5_ ( .J(n43), .K(n43), .TI(shifter_N11), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(shifter_temp_5_) );
  GTECH_FJK2S shifter_temp_reg_4_ ( .J(n43), .K(n43), .TI(shifter_N10), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(shifter_temp_4_) );
  GTECH_FJK2S shifter_temp_reg_3_ ( .J(n43), .K(n43), .TI(shifter_N9), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(shifter_temp_3_) );
  GTECH_FJK2S shifter_temp_reg_2_ ( .J(n43), .K(n43), .TI(shifter_N8), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(shifter_temp_2_) );
  GTECH_FJK2S shifter_temp_reg_1_ ( .J(n43), .K(n43), .TI(shifter_N7), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(shifter_temp_1_) );
  GTECH_FJK2S shifter_temp_reg_0_ ( .J(n43), .K(n43), .TI(shifter_N6), .TE(
        shifter_N22), .CP(clk), .CD(n132), .Q(lsb), .QN(n137) );
  GTECH_FJK2S controller_out_cmd_reg ( .J(n43), .K(n43), .TI(controller_N92), 
        .TE(controller_N95), .CP(clk), .CD(n132), .Q(out_cmd) );
  GTECH_ZERO U157 ( .Z(n43) );
  GTECH_ONE U158 ( .Z(n127) );
  GTECH_OAI2N2 U159 ( .A(n172), .B(n173), .C(Q[3]), .D(n174), .Z(shifter_N9)
         );
  GTECH_NOT U160 ( .A(shifter_temp_4_), .Z(n173) );
  GTECH_OAI2N2 U161 ( .A(n172), .B(n175), .C(Q[2]), .D(n174), .Z(shifter_N8)
         );
  GTECH_NOT U162 ( .A(shifter_temp_3_), .Z(n175) );
  GTECH_OAI2N2 U163 ( .A(n172), .B(n176), .C(Q[1]), .D(n174), .Z(shifter_N7)
         );
  GTECH_NOT U164 ( .A(shifter_temp_2_), .Z(n176) );
  GTECH_OAI2N2 U165 ( .A(n172), .B(n177), .C(Q[0]), .D(n174), .Z(shifter_N6)
         );
  GTECH_NOT U166 ( .A(shifter_temp_1_), .Z(n177) );
  GTECH_NOT U167 ( .A(n178), .Z(shifter_N24) );
  GTECH_NAND2 U168 ( .A(n178), .B(n179), .Z(shifter_N23) );
  GTECH_NAND2 U169 ( .A(n136), .B(n180), .Z(n178) );
  GTECH_NOT U170 ( .A(n135), .Z(n180) );
  GTECH_NAND2 U171 ( .A(n172), .B(n136), .Z(shifter_N22) );
  GTECH_AND2 U172 ( .A(n181), .B(n182), .Z(shifter_N21) );
  GTECH_OAI22 U173 ( .A(n183), .B(n184), .C(n12), .D(n185), .Z(n182) );
  GTECH_NOT U174 ( .A(n179), .Z(n181) );
  GTECH_OAI22 U175 ( .A(n12), .B(n186), .C(n187), .D(n179), .Z(shifter_N20) );
  GTECH_AOI222 U176 ( .A(n185), .B(n188), .C(n189), .D(n183), .E(n190), .F(
        n191), .Z(n187) );
  GTECH_XOR2 U177 ( .A(n12), .B(D[7]), .Z(n190) );
  GTECH_AND2 U178 ( .A(n12), .B(D[7]), .Z(n189) );
  GTECH_NOT U179 ( .A(n192), .Z(n185) );
  GTECH_NAND2 U180 ( .A(n183), .B(n184), .Z(n192) );
  GTECH_NOT U181 ( .A(D[7]), .Z(n184) );
  GTECH_NOT U182 ( .A(n191), .Z(n183) );
  GTECH_OAI21 U183 ( .A(n13), .B(n193), .C(n194), .Z(n191) );
  GTECH_OAI21 U184 ( .A(D[6]), .B(n195), .C(n196), .Z(n194) );
  GTECH_NOT U185 ( .A(D[6]), .Z(n193) );
  GTECH_OAI22 U186 ( .A(n13), .B(n186), .C(n197), .D(n179), .Z(shifter_N19) );
  GTECH_XOR3 U187 ( .A(n13), .B(D[6]), .C(n196), .Z(n197) );
  GTECH_OAI21 U188 ( .A(n14), .B(n198), .C(n199), .Z(n196) );
  GTECH_OAI21 U189 ( .A(D[5]), .B(n200), .C(n201), .Z(n199) );
  GTECH_NOT U190 ( .A(D[5]), .Z(n198) );
  GTECH_OAI22 U191 ( .A(n14), .B(n186), .C(n202), .D(n179), .Z(shifter_N18) );
  GTECH_XOR3 U192 ( .A(n14), .B(D[5]), .C(n201), .Z(n202) );
  GTECH_OAI21 U193 ( .A(n15), .B(n203), .C(n204), .Z(n201) );
  GTECH_OAI21 U194 ( .A(D[4]), .B(n205), .C(n206), .Z(n204) );
  GTECH_NOT U195 ( .A(D[4]), .Z(n203) );
  GTECH_OAI22 U196 ( .A(n15), .B(n186), .C(n207), .D(n179), .Z(shifter_N17) );
  GTECH_XOR3 U197 ( .A(n15), .B(D[4]), .C(n206), .Z(n207) );
  GTECH_OAI21 U198 ( .A(n16), .B(n208), .C(n209), .Z(n206) );
  GTECH_OAI21 U199 ( .A(D[3]), .B(n210), .C(n211), .Z(n209) );
  GTECH_NOT U200 ( .A(D[3]), .Z(n208) );
  GTECH_OAI22 U201 ( .A(n16), .B(n186), .C(n212), .D(n179), .Z(shifter_N16) );
  GTECH_XOR3 U202 ( .A(n16), .B(D[3]), .C(n211), .Z(n212) );
  GTECH_OAI21 U203 ( .A(n17), .B(n213), .C(n214), .Z(n211) );
  GTECH_OAI21 U204 ( .A(D[2]), .B(n215), .C(n216), .Z(n214) );
  GTECH_NOT U205 ( .A(D[2]), .Z(n213) );
  GTECH_OAI22 U206 ( .A(n17), .B(n186), .C(n217), .D(n179), .Z(shifter_N15) );
  GTECH_XOR3 U207 ( .A(n17), .B(D[2]), .C(n216), .Z(n217) );
  GTECH_OAI21 U208 ( .A(n18), .B(n218), .C(n219), .Z(n216) );
  GTECH_OAI21 U209 ( .A(D[1]), .B(n220), .C(n221), .Z(n219) );
  GTECH_NOT U210 ( .A(D[1]), .Z(n218) );
  GTECH_OAI22 U211 ( .A(n18), .B(n186), .C(n179), .D(n222), .Z(shifter_N14) );
  GTECH_XOR3 U212 ( .A(n18), .B(D[1]), .C(n221), .Z(n222) );
  GTECH_NOT U213 ( .A(n223), .Z(n221) );
  GTECH_NAND2 U214 ( .A(D[0]), .B(n224), .Z(n223) );
  GTECH_AO21 U215 ( .A(Q[7]), .B(n174), .C(n225), .Z(shifter_N13) );
  GTECH_OAI22 U216 ( .A(n179), .B(n226), .C(n11), .D(n186), .Z(n225) );
  GTECH_XOR2 U217 ( .A(D[0]), .B(n11), .Z(n226) );
  GTECH_OAI2N2 U218 ( .A(n172), .B(n227), .C(Q[6]), .D(n174), .Z(shifter_N12)
         );
  GTECH_NOT U219 ( .A(shifter_temp_7_), .Z(n227) );
  GTECH_OAI2N2 U220 ( .A(n172), .B(n228), .C(Q[5]), .D(n174), .Z(shifter_N11)
         );
  GTECH_NOT U221 ( .A(shifter_temp_6_), .Z(n228) );
  GTECH_OAI2N2 U222 ( .A(n172), .B(n229), .C(Q[4]), .D(n174), .Z(shifter_N10)
         );
  GTECH_NOT U223 ( .A(n136), .Z(n174) );
  GTECH_NOT U224 ( .A(shifter_temp_5_), .Z(n229) );
  GTECH_NOT U225 ( .A(n230), .Z(n172) );
  GTECH_NAND2 U226 ( .A(n186), .B(n179), .Z(n230) );
  GTECH_NAND4 U227 ( .A(shifter_add_temp), .B(shift_cmd), .C(n136), .D(n135), 
        .Z(n179) );
  GTECH_NAND4 U228 ( .A(shift_cmd), .B(n136), .C(n135), .D(n231), .Z(n186) );
  GTECH_NOT U229 ( .A(shifter_add_temp), .Z(n231) );
  GTECH_AND2 U230 ( .A(out_cmd), .B(n220), .Z(out[9]) );
  GTECH_NOT U231 ( .A(n18), .Z(n220) );
  GTECH_AND2 U232 ( .A(out_cmd), .B(n224), .Z(out[8]) );
  GTECH_NOT U233 ( .A(n11), .Z(n224) );
  GTECH_AND2 U234 ( .A(out_cmd), .B(shifter_temp_7_), .Z(out[7]) );
  GTECH_AND2 U235 ( .A(out_cmd), .B(shifter_temp_6_), .Z(out[6]) );
  GTECH_AND2 U236 ( .A(out_cmd), .B(shifter_temp_5_), .Z(out[5]) );
  GTECH_AND2 U237 ( .A(out_cmd), .B(shifter_temp_4_), .Z(out[4]) );
  GTECH_AND2 U238 ( .A(out_cmd), .B(shifter_temp_3_), .Z(out[3]) );
  GTECH_AND2 U239 ( .A(out_cmd), .B(shifter_temp_2_), .Z(out[2]) );
  GTECH_AND2 U240 ( .A(out_cmd), .B(shifter_temp_1_), .Z(out[1]) );
  GTECH_AND2 U241 ( .A(out_cmd), .B(n188), .Z(out[15]) );
  GTECH_NOT U242 ( .A(n12), .Z(n188) );
  GTECH_AND2 U243 ( .A(out_cmd), .B(n195), .Z(out[14]) );
  GTECH_NOT U244 ( .A(n13), .Z(n195) );
  GTECH_AND2 U245 ( .A(out_cmd), .B(n200), .Z(out[13]) );
  GTECH_NOT U246 ( .A(n14), .Z(n200) );
  GTECH_AND2 U247 ( .A(out_cmd), .B(n205), .Z(out[12]) );
  GTECH_NOT U248 ( .A(n15), .Z(n205) );
  GTECH_AND2 U249 ( .A(out_cmd), .B(n210), .Z(out[11]) );
  GTECH_NOT U250 ( .A(n16), .Z(n210) );
  GTECH_AND2 U251 ( .A(out_cmd), .B(n215), .Z(out[10]) );
  GTECH_NOT U252 ( .A(n17), .Z(n215) );
  GTECH_AND2 U253 ( .A(out_cmd), .B(n232), .Z(out[0]) );
  GTECH_AND2 U254 ( .A(controller_N98), .B(n233), .Z(controller_N97) );
  GTECH_NOT U255 ( .A(n234), .Z(controller_N98) );
  GTECH_OAI21 U256 ( .A(n235), .B(n232), .C(n236), .Z(controller_N96) );
  GTECH_OAI21 U257 ( .A(n233), .B(n234), .C(n237), .Z(controller_N94) );
  GTECH_AND2 U258 ( .A(n238), .B(n239), .Z(n237) );
  GTECH_NAND3 U259 ( .A(n138), .B(n232), .C(n240), .Z(n238) );
  GTECH_AND3 U260 ( .A(n138), .B(n241), .C(n139), .Z(controller_N93) );
  GTECH_AOI2N2 U261 ( .A(n8), .B(n129), .C(n232), .D(n8), .Z(n241) );
  GTECH_NOT U262 ( .A(n137), .Z(n232) );
  GTECH_AND4 U263 ( .A(n129), .B(n139), .C(n8), .D(n138), .Z(controller_N92)
         );
  GTECH_NOT U264 ( .A(n236), .Z(controller_N91) );
  GTECH_NAND2 U265 ( .A(n240), .B(n242), .Z(n236) );
  GTECH_NOT U266 ( .A(n235), .Z(n240) );
  GTECH_NAND2 U267 ( .A(n139), .B(n243), .Z(n235) );
  GTECH_NOT U268 ( .A(n8), .Z(n243) );
  GTECH_NOT U269 ( .A(n239), .Z(controller_N90) );
  GTECH_NAND3 U270 ( .A(n8), .B(n242), .C(n139), .Z(n239) );
  GTECH_NOT U271 ( .A(n138), .Z(n242) );
  GTECH_AOI21 U272 ( .A(n244), .B(n245), .C(n153), .Z(controller_N83) );
  GTECH_NOT U273 ( .A(n152), .Z(n245) );
  GTECH_NOT U274 ( .A(n246), .Z(n244) );
  GTECH_AND2 U275 ( .A(n247), .B(n248), .Z(controller_N82) );
  GTECH_XOR2 U276 ( .A(n246), .B(n152), .Z(n247) );
  GTECH_NAND2 U277 ( .A(n249), .B(n250), .Z(n246) );
  GTECH_NOT U278 ( .A(n151), .Z(n250) );
  GTECH_NOT U279 ( .A(n251), .Z(n249) );
  GTECH_AND2 U280 ( .A(n252), .B(n248), .Z(controller_N81) );
  GTECH_XOR2 U281 ( .A(n251), .B(n151), .Z(n252) );
  GTECH_NAND2 U282 ( .A(n253), .B(n254), .Z(n251) );
  GTECH_NOT U283 ( .A(n150), .Z(n254) );
  GTECH_NOT U284 ( .A(n255), .Z(n253) );
  GTECH_AND2 U285 ( .A(n256), .B(n248), .Z(controller_N80) );
  GTECH_XOR2 U286 ( .A(n255), .B(n150), .Z(n256) );
  GTECH_NAND2 U287 ( .A(n257), .B(n258), .Z(n255) );
  GTECH_NOT U288 ( .A(n149), .Z(n258) );
  GTECH_NOT U289 ( .A(n259), .Z(n257) );
  GTECH_AND2 U290 ( .A(n260), .B(n248), .Z(controller_N79) );
  GTECH_XOR2 U291 ( .A(n259), .B(n149), .Z(n260) );
  GTECH_NAND2 U292 ( .A(n261), .B(n262), .Z(n259) );
  GTECH_NOT U293 ( .A(n148), .Z(n262) );
  GTECH_NOT U294 ( .A(n263), .Z(n261) );
  GTECH_AND2 U295 ( .A(n264), .B(n248), .Z(controller_N78) );
  GTECH_XOR2 U296 ( .A(n263), .B(n148), .Z(n264) );
  GTECH_NAND2 U297 ( .A(n265), .B(n266), .Z(n263) );
  GTECH_NOT U298 ( .A(n147), .Z(n266) );
  GTECH_NOT U299 ( .A(n267), .Z(n265) );
  GTECH_AND2 U300 ( .A(n268), .B(n248), .Z(controller_N77) );
  GTECH_XOR2 U301 ( .A(n267), .B(n147), .Z(n268) );
  GTECH_NAND2 U302 ( .A(n269), .B(n270), .Z(n267) );
  GTECH_NOT U303 ( .A(n146), .Z(n270) );
  GTECH_NOT U304 ( .A(n271), .Z(n269) );
  GTECH_AND2 U305 ( .A(n272), .B(n248), .Z(controller_N76) );
  GTECH_XOR2 U306 ( .A(n271), .B(n146), .Z(n272) );
  GTECH_NAND2 U307 ( .A(n273), .B(n274), .Z(n271) );
  GTECH_NOT U308 ( .A(n145), .Z(n274) );
  GTECH_NOT U309 ( .A(n275), .Z(n273) );
  GTECH_AND2 U310 ( .A(n276), .B(n248), .Z(controller_N75) );
  GTECH_XOR2 U311 ( .A(n275), .B(n145), .Z(n276) );
  GTECH_NAND2 U312 ( .A(n277), .B(n278), .Z(n275) );
  GTECH_NOT U313 ( .A(n144), .Z(n278) );
  GTECH_NOT U314 ( .A(n279), .Z(n277) );
  GTECH_AND2 U315 ( .A(n280), .B(n248), .Z(controller_N74) );
  GTECH_XOR2 U316 ( .A(n279), .B(n144), .Z(n280) );
  GTECH_NAND2 U317 ( .A(n281), .B(n282), .Z(n279) );
  GTECH_NOT U318 ( .A(n143), .Z(n282) );
  GTECH_NOT U319 ( .A(n283), .Z(n281) );
  GTECH_AND2 U320 ( .A(n284), .B(n248), .Z(controller_N73) );
  GTECH_XOR2 U321 ( .A(n283), .B(n143), .Z(n284) );
  GTECH_NAND2 U322 ( .A(n285), .B(n286), .Z(n283) );
  GTECH_NOT U323 ( .A(n142), .Z(n286) );
  GTECH_NOT U324 ( .A(n287), .Z(n285) );
  GTECH_AND2 U325 ( .A(n288), .B(n248), .Z(controller_N72) );
  GTECH_XOR2 U326 ( .A(n287), .B(n142), .Z(n288) );
  GTECH_NAND2 U327 ( .A(n289), .B(n290), .Z(n287) );
  GTECH_NOT U328 ( .A(n141), .Z(n290) );
  GTECH_NOT U329 ( .A(n291), .Z(n289) );
  GTECH_AND2 U330 ( .A(n292), .B(n248), .Z(controller_N71) );
  GTECH_XOR2 U331 ( .A(n291), .B(n141), .Z(n292) );
  GTECH_NAND2 U332 ( .A(n293), .B(n294), .Z(n291) );
  GTECH_NOT U333 ( .A(n140), .Z(n294) );
  GTECH_NOT U334 ( .A(n295), .Z(n293) );
  GTECH_AND2 U335 ( .A(n296), .B(n248), .Z(controller_N70) );
  GTECH_XOR2 U336 ( .A(n295), .B(n140), .Z(n296) );
  GTECH_NAND2 U337 ( .A(n297), .B(n298), .Z(n295) );
  GTECH_NOT U338 ( .A(n171), .Z(n298) );
  GTECH_NOT U339 ( .A(n299), .Z(n297) );
  GTECH_AND2 U340 ( .A(n300), .B(n248), .Z(controller_N69) );
  GTECH_XOR2 U341 ( .A(n299), .B(n171), .Z(n300) );
  GTECH_NAND2 U342 ( .A(n301), .B(n302), .Z(n299) );
  GTECH_NOT U343 ( .A(n170), .Z(n302) );
  GTECH_NOT U344 ( .A(n303), .Z(n301) );
  GTECH_AND2 U345 ( .A(n304), .B(n248), .Z(controller_N68) );
  GTECH_XOR2 U346 ( .A(n303), .B(n170), .Z(n304) );
  GTECH_NAND2 U347 ( .A(n305), .B(n306), .Z(n303) );
  GTECH_NOT U348 ( .A(n169), .Z(n306) );
  GTECH_NOT U349 ( .A(n307), .Z(n305) );
  GTECH_AND2 U350 ( .A(n308), .B(n248), .Z(controller_N67) );
  GTECH_XOR2 U351 ( .A(n307), .B(n169), .Z(n308) );
  GTECH_NAND2 U352 ( .A(n309), .B(n310), .Z(n307) );
  GTECH_NOT U353 ( .A(n168), .Z(n310) );
  GTECH_NOT U354 ( .A(n311), .Z(n309) );
  GTECH_AND2 U355 ( .A(n312), .B(n248), .Z(controller_N66) );
  GTECH_XOR2 U356 ( .A(n311), .B(n168), .Z(n312) );
  GTECH_NAND2 U357 ( .A(n313), .B(n314), .Z(n311) );
  GTECH_NOT U358 ( .A(n167), .Z(n314) );
  GTECH_NOT U359 ( .A(n315), .Z(n313) );
  GTECH_AND2 U360 ( .A(n316), .B(n248), .Z(controller_N65) );
  GTECH_XOR2 U361 ( .A(n315), .B(n167), .Z(n316) );
  GTECH_NAND2 U362 ( .A(n317), .B(n318), .Z(n315) );
  GTECH_NOT U363 ( .A(n166), .Z(n318) );
  GTECH_NOT U364 ( .A(n319), .Z(n317) );
  GTECH_AND2 U365 ( .A(n320), .B(n248), .Z(controller_N64) );
  GTECH_XOR2 U366 ( .A(n319), .B(n166), .Z(n320) );
  GTECH_NAND2 U367 ( .A(n321), .B(n322), .Z(n319) );
  GTECH_NOT U368 ( .A(n165), .Z(n322) );
  GTECH_NOT U369 ( .A(n323), .Z(n321) );
  GTECH_AND2 U370 ( .A(n324), .B(n248), .Z(controller_N63) );
  GTECH_XOR2 U371 ( .A(n323), .B(n165), .Z(n324) );
  GTECH_NAND2 U372 ( .A(n325), .B(n326), .Z(n323) );
  GTECH_NOT U373 ( .A(n164), .Z(n326) );
  GTECH_NOT U374 ( .A(n327), .Z(n325) );
  GTECH_AND2 U375 ( .A(n328), .B(n248), .Z(controller_N62) );
  GTECH_XOR2 U376 ( .A(n327), .B(n164), .Z(n328) );
  GTECH_NAND2 U377 ( .A(n329), .B(n330), .Z(n327) );
  GTECH_NOT U378 ( .A(n163), .Z(n330) );
  GTECH_NOT U379 ( .A(n331), .Z(n329) );
  GTECH_AND2 U380 ( .A(n332), .B(n248), .Z(controller_N61) );
  GTECH_XOR2 U381 ( .A(n331), .B(n163), .Z(n332) );
  GTECH_NAND2 U382 ( .A(n333), .B(n334), .Z(n331) );
  GTECH_NOT U383 ( .A(n162), .Z(n334) );
  GTECH_NOT U384 ( .A(n335), .Z(n333) );
  GTECH_AND2 U385 ( .A(n336), .B(n248), .Z(controller_N60) );
  GTECH_XOR2 U386 ( .A(n335), .B(n162), .Z(n336) );
  GTECH_NAND2 U387 ( .A(n337), .B(n338), .Z(n335) );
  GTECH_NOT U388 ( .A(n161), .Z(n338) );
  GTECH_NOT U389 ( .A(n339), .Z(n337) );
  GTECH_AND2 U390 ( .A(n340), .B(n248), .Z(controller_N59) );
  GTECH_XOR2 U391 ( .A(n339), .B(n161), .Z(n340) );
  GTECH_NAND2 U392 ( .A(n341), .B(n342), .Z(n339) );
  GTECH_NOT U393 ( .A(n160), .Z(n342) );
  GTECH_NOT U394 ( .A(n343), .Z(n341) );
  GTECH_AND2 U395 ( .A(n344), .B(n248), .Z(controller_N58) );
  GTECH_XOR2 U396 ( .A(n343), .B(n160), .Z(n344) );
  GTECH_NAND2 U397 ( .A(n345), .B(n346), .Z(n343) );
  GTECH_NOT U398 ( .A(n159), .Z(n346) );
  GTECH_NOT U399 ( .A(n347), .Z(n345) );
  GTECH_AND2 U400 ( .A(n348), .B(n248), .Z(controller_N57) );
  GTECH_XOR2 U401 ( .A(n347), .B(n159), .Z(n348) );
  GTECH_NAND2 U402 ( .A(n349), .B(n350), .Z(n347) );
  GTECH_NOT U403 ( .A(n158), .Z(n350) );
  GTECH_NOT U404 ( .A(n351), .Z(n349) );
  GTECH_AND2 U405 ( .A(n352), .B(n248), .Z(controller_N56) );
  GTECH_XOR2 U406 ( .A(n351), .B(n158), .Z(n352) );
  GTECH_NAND2 U407 ( .A(n353), .B(n354), .Z(n351) );
  GTECH_NOT U408 ( .A(n157), .Z(n354) );
  GTECH_NOT U409 ( .A(n355), .Z(n353) );
  GTECH_AND2 U410 ( .A(n356), .B(n248), .Z(controller_N55) );
  GTECH_XOR2 U411 ( .A(n355), .B(n157), .Z(n356) );
  GTECH_NAND3 U412 ( .A(n357), .B(n358), .C(n359), .Z(n355) );
  GTECH_NOT U413 ( .A(n156), .Z(n358) );
  GTECH_NOT U414 ( .A(n155), .Z(n357) );
  GTECH_OAI22 U415 ( .A(n156), .B(n360), .C(n233), .D(n361), .Z(controller_N54) );
  GTECH_OAI21 U416 ( .A(n156), .B(n155), .C(n362), .Z(n361) );
  GTECH_OAI21 U417 ( .A(n155), .B(n154), .C(n156), .Z(n362) );
  GTECH_NOT U418 ( .A(n248), .Z(n233) );
  GTECH_OAI21 U419 ( .A(n155), .B(n360), .C(n363), .Z(controller_N53) );
  GTECH_NAND3 U420 ( .A(n248), .B(n359), .C(n155), .Z(n363) );
  GTECH_NOT U421 ( .A(n154), .Z(n359) );
  GTECH_NOT U422 ( .A(n360), .Z(controller_N52) );
  GTECH_NAND2 U423 ( .A(n154), .B(n248), .Z(n360) );
  GTECH_OAI21 U424 ( .A(n364), .B(n365), .C(n153), .Z(n248) );
  GTECH_NAND8 U425 ( .A(n170), .B(n169), .C(n171), .D(n366), .E(n163), .F(n162), .G(n164), .H(n367), .Z(n365) );
  GTECH_AND4 U426 ( .A(n161), .B(n160), .C(n159), .D(n158), .Z(n367) );
  GTECH_AND4 U427 ( .A(n168), .B(n167), .C(n166), .D(n165), .Z(n366) );
  GTECH_NAND8 U428 ( .A(n152), .B(n151), .C(n157), .D(n368), .E(n145), .F(n144), .G(n146), .H(n369), .Z(n364) );
  GTECH_AND4 U429 ( .A(n143), .B(n142), .C(n141), .D(n140), .Z(n369) );
  GTECH_AND4 U430 ( .A(n150), .B(n149), .C(n148), .D(n147), .Z(n368) );
  GTECH_AND2 U431 ( .A(controller_N95), .B(n132), .Z(controller_N102) );
  GTECH_NOT U432 ( .A(rst), .Z(n132) );
  GTECH_NAND2 U433 ( .A(n370), .B(n234), .Z(controller_N95) );
  GTECH_NAND3 U434 ( .A(n138), .B(n370), .C(n8), .Z(n234) );
  GTECH_NOT U435 ( .A(n139), .Z(n370) );
endmodule

