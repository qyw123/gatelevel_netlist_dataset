
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374;

  GTECH_MUX2 U132 ( .A(n271), .B(n272), .S(n273), .Z(sum[9]) );
  GTECH_XNOR2 U133 ( .A(n274), .B(n275), .Z(n272) );
  GTECH_XNOR2 U134 ( .A(n276), .B(n275), .Z(n271) );
  GTECH_OA21 U135 ( .A(b[9]), .B(a[9]), .C(n277), .Z(n275) );
  GTECH_XNOR2 U136 ( .A(n278), .B(n273), .Z(sum[8]) );
  GTECH_MUX2 U137 ( .A(n279), .B(n280), .S(n281), .Z(sum[7]) );
  GTECH_XNOR2 U138 ( .A(n282), .B(n283), .Z(n280) );
  GTECH_OA21 U139 ( .A(n284), .B(n285), .C(n286), .Z(n283) );
  GTECH_XNOR2 U140 ( .A(n282), .B(n287), .Z(n279) );
  GTECH_XOR2 U141 ( .A(a[7]), .B(b[7]), .Z(n282) );
  GTECH_MUX2 U142 ( .A(n288), .B(n289), .S(n281), .Z(sum[6]) );
  GTECH_XNOR2 U143 ( .A(n290), .B(n285), .Z(n289) );
  GTECH_AO21 U144 ( .A(n291), .B(n292), .C(n293), .Z(n285) );
  GTECH_XNOR2 U145 ( .A(n290), .B(n294), .Z(n288) );
  GTECH_AND_NOT U146 ( .A(n286), .B(n284), .Z(n290) );
  GTECH_MUX2 U147 ( .A(n295), .B(n296), .S(n281), .Z(sum[5]) );
  GTECH_XNOR2 U148 ( .A(n291), .B(n297), .Z(n296) );
  GTECH_XOR2 U149 ( .A(n298), .B(n297), .Z(n295) );
  GTECH_OA21 U150 ( .A(b[5]), .B(a[5]), .C(n292), .Z(n297) );
  GTECH_OR_NOT U151 ( .A(n299), .B(n300), .Z(sum[4]) );
  GTECH_AO21 U152 ( .A(n298), .B(n291), .C(n281), .Z(n300) );
  GTECH_MUX2 U153 ( .A(n301), .B(n302), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U154 ( .A(n303), .B(n304), .Z(n302) );
  GTECH_XOR2 U155 ( .A(n303), .B(n305), .Z(n301) );
  GTECH_AOI21 U156 ( .A(n306), .B(n307), .C(n308), .Z(n305) );
  GTECH_XNOR2 U157 ( .A(a[3]), .B(b[3]), .Z(n303) );
  GTECH_MUX2 U158 ( .A(n309), .B(n310), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U159 ( .A(n311), .B(n312), .Z(n310) );
  GTECH_XOR2 U160 ( .A(n311), .B(n307), .Z(n309) );
  GTECH_OA21 U161 ( .A(n313), .B(n314), .C(n315), .Z(n307) );
  GTECH_AND_NOT U162 ( .A(n306), .B(n308), .Z(n311) );
  GTECH_MUX2 U163 ( .A(n316), .B(n317), .S(n318), .Z(sum[1]) );
  GTECH_OA21 U164 ( .A(a[1]), .B(b[1]), .C(n319), .Z(n318) );
  GTECH_NOT U165 ( .A(n314), .Z(n319) );
  GTECH_NOT U166 ( .A(n320), .Z(n317) );
  GTECH_OA21 U167 ( .A(n313), .B(cin), .C(n321), .Z(n320) );
  GTECH_AO21 U168 ( .A(cin), .B(n321), .C(n313), .Z(n316) );
  GTECH_AND2 U169 ( .A(a[0]), .B(b[0]), .Z(n313) );
  GTECH_MUX2 U170 ( .A(n322), .B(n323), .S(n324), .Z(sum[15]) );
  GTECH_XOR2 U171 ( .A(n325), .B(n326), .Z(n323) );
  GTECH_XOR2 U172 ( .A(n325), .B(n327), .Z(n322) );
  GTECH_OA21 U173 ( .A(n328), .B(n329), .C(n330), .Z(n327) );
  GTECH_XNOR2 U174 ( .A(n331), .B(n332), .Z(n325) );
  GTECH_MUX2 U175 ( .A(n333), .B(n334), .S(n324), .Z(sum[14]) );
  GTECH_XNOR2 U176 ( .A(n335), .B(n336), .Z(n334) );
  GTECH_XNOR2 U177 ( .A(n335), .B(n329), .Z(n333) );
  GTECH_AO21 U178 ( .A(n337), .B(n338), .C(n339), .Z(n329) );
  GTECH_AND_NOT U179 ( .A(n330), .B(n328), .Z(n335) );
  GTECH_MUX2 U180 ( .A(n340), .B(n341), .S(n324), .Z(sum[13]) );
  GTECH_XOR2 U181 ( .A(n342), .B(n343), .Z(n341) );
  GTECH_XNOR2 U182 ( .A(n342), .B(n337), .Z(n340) );
  GTECH_OA21 U183 ( .A(b[13]), .B(a[13]), .C(n338), .Z(n342) );
  GTECH_OR_NOT U184 ( .A(n344), .B(n345), .Z(sum[12]) );
  GTECH_AO21 U185 ( .A(n343), .B(n337), .C(n346), .Z(n345) );
  GTECH_MUX2 U186 ( .A(n347), .B(n348), .S(n273), .Z(sum[11]) );
  GTECH_XOR2 U187 ( .A(n349), .B(n350), .Z(n348) );
  GTECH_OA21 U188 ( .A(n351), .B(n352), .C(n353), .Z(n350) );
  GTECH_XOR2 U189 ( .A(n349), .B(n354), .Z(n347) );
  GTECH_XNOR2 U190 ( .A(a[11]), .B(b[11]), .Z(n349) );
  GTECH_MUX2 U191 ( .A(n355), .B(n356), .S(n273), .Z(sum[10]) );
  GTECH_XNOR2 U192 ( .A(n357), .B(n352), .Z(n356) );
  GTECH_AO21 U193 ( .A(n274), .B(n277), .C(n358), .Z(n352) );
  GTECH_XNOR2 U194 ( .A(n357), .B(n359), .Z(n355) );
  GTECH_AND_NOT U195 ( .A(n353), .B(n351), .Z(n357) );
  GTECH_XNOR2 U196 ( .A(cin), .B(n360), .Z(sum[0]) );
  GTECH_AO21 U197 ( .A(n324), .B(n361), .C(n344), .Z(cout) );
  GTECH_AND3 U198 ( .A(n337), .B(n343), .C(n346), .Z(n344) );
  GTECH_NOT U199 ( .A(n324), .Z(n346) );
  GTECH_NOT U200 ( .A(n362), .Z(n343) );
  GTECH_NAND2 U201 ( .A(a[12]), .B(b[12]), .Z(n337) );
  GTECH_OAI22 U202 ( .A(n326), .B(n331), .C(n363), .D(n332), .Z(n361) );
  GTECH_NOT U203 ( .A(b[15]), .Z(n332) );
  GTECH_AND_NOT U204 ( .A(n326), .B(a[15]), .Z(n363) );
  GTECH_NOT U205 ( .A(a[15]), .Z(n331) );
  GTECH_OA21 U206 ( .A(n336), .B(n328), .C(n330), .Z(n326) );
  GTECH_NAND2 U207 ( .A(b[14]), .B(a[14]), .Z(n330) );
  GTECH_NOR2 U208 ( .A(a[14]), .B(b[14]), .Z(n328) );
  GTECH_AO21 U209 ( .A(n362), .B(n338), .C(n339), .Z(n336) );
  GTECH_NOR2 U210 ( .A(a[13]), .B(b[13]), .Z(n339) );
  GTECH_NAND2 U211 ( .A(b[13]), .B(a[13]), .Z(n338) );
  GTECH_NOR2 U212 ( .A(b[12]), .B(a[12]), .Z(n362) );
  GTECH_MUX2 U213 ( .A(n364), .B(n278), .S(n273), .Z(n324) );
  GTECH_AOI21 U214 ( .A(n365), .B(n366), .C(n299), .Z(n273) );
  GTECH_AND3 U215 ( .A(n298), .B(n291), .C(n281), .Z(n299) );
  GTECH_NAND2 U216 ( .A(b[4]), .B(a[4]), .Z(n291) );
  GTECH_NOT U217 ( .A(n367), .Z(n298) );
  GTECH_OAI2N2 U218 ( .A(n287), .B(n368), .C(n369), .D(b[7]), .Z(n366) );
  GTECH_OR_NOT U219 ( .A(a[7]), .B(n287), .Z(n369) );
  GTECH_NOT U220 ( .A(a[7]), .Z(n368) );
  GTECH_OA21 U221 ( .A(n294), .B(n284), .C(n286), .Z(n287) );
  GTECH_NAND2 U222 ( .A(b[6]), .B(a[6]), .Z(n286) );
  GTECH_NOR2 U223 ( .A(a[6]), .B(b[6]), .Z(n284) );
  GTECH_AO21 U224 ( .A(n367), .B(n292), .C(n293), .Z(n294) );
  GTECH_NOR2 U225 ( .A(b[5]), .B(a[5]), .Z(n293) );
  GTECH_NAND2 U226 ( .A(a[5]), .B(b[5]), .Z(n292) );
  GTECH_NOR2 U227 ( .A(a[4]), .B(b[4]), .Z(n367) );
  GTECH_NOT U228 ( .A(n281), .Z(n365) );
  GTECH_MUX2 U229 ( .A(n360), .B(n370), .S(cin), .Z(n281) );
  GTECH_AOI21 U230 ( .A(n304), .B(a[3]), .C(n371), .Z(n370) );
  GTECH_OA21 U231 ( .A(n304), .B(a[3]), .C(b[3]), .Z(n371) );
  GTECH_AO21 U232 ( .A(n312), .B(n306), .C(n308), .Z(n304) );
  GTECH_AND2 U233 ( .A(b[2]), .B(a[2]), .Z(n308) );
  GTECH_OR2 U234 ( .A(a[2]), .B(b[2]), .Z(n306) );
  GTECH_OA21 U235 ( .A(n321), .B(n314), .C(n315), .Z(n312) );
  GTECH_OR2 U236 ( .A(a[1]), .B(b[1]), .Z(n315) );
  GTECH_AND2 U237 ( .A(b[1]), .B(a[1]), .Z(n314) );
  GTECH_OR2 U238 ( .A(a[0]), .B(b[0]), .Z(n321) );
  GTECH_XOR2 U239 ( .A(a[0]), .B(n372), .Z(n360) );
  GTECH_NOT U240 ( .A(b[0]), .Z(n372) );
  GTECH_AND_NOT U241 ( .A(n274), .B(n276), .Z(n278) );
  GTECH_NAND2 U242 ( .A(a[8]), .B(b[8]), .Z(n274) );
  GTECH_OA21 U243 ( .A(a[11]), .B(n373), .C(n374), .Z(n364) );
  GTECH_AO21 U244 ( .A(a[11]), .B(n373), .C(b[11]), .Z(n374) );
  GTECH_NOT U245 ( .A(n354), .Z(n373) );
  GTECH_OA21 U246 ( .A(n359), .B(n351), .C(n353), .Z(n354) );
  GTECH_NAND2 U247 ( .A(b[10]), .B(a[10]), .Z(n353) );
  GTECH_NOR2 U248 ( .A(a[10]), .B(b[10]), .Z(n351) );
  GTECH_AO21 U249 ( .A(n276), .B(n277), .C(n358), .Z(n359) );
  GTECH_NOR2 U250 ( .A(b[9]), .B(a[9]), .Z(n358) );
  GTECH_NAND2 U251 ( .A(a[9]), .B(b[9]), .Z(n277) );
  GTECH_NOR2 U252 ( .A(b[8]), .B(a[8]), .Z(n276) );
endmodule

