
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n128, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n128), .K(n128), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n265) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n128), .K(n128), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n128), .K(n128), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n128), .K(n128), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n128), .K(n128), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n128), .K(n128), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]), .QN(n282) );
  GTECH_FJK1S A_reg_15_ ( .J(n128), .K(n128), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n281) );
  GTECH_FJK1S A_reg_14_ ( .J(n128), .K(n128), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n280) );
  GTECH_FJK1S A_reg_13_ ( .J(n128), .K(n128), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n279) );
  GTECH_FJK1S A_reg_12_ ( .J(n128), .K(n128), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n278) );
  GTECH_FJK1S A_reg_11_ ( .J(n128), .K(n128), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n277) );
  GTECH_FJK1S A_reg_10_ ( .J(n128), .K(n128), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n276) );
  GTECH_FJK1S A_reg_9_ ( .J(n128), .K(n128), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n275) );
  GTECH_FJK1S A_reg_8_ ( .J(n128), .K(n128), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n274) );
  GTECH_FJK1S A_reg_7_ ( .J(n128), .K(n128), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n273) );
  GTECH_FJK1S A_reg_6_ ( .J(n128), .K(n128), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n272) );
  GTECH_FJK1S A_reg_5_ ( .J(n128), .K(n128), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n271) );
  GTECH_FJK1S A_reg_4_ ( .J(n128), .K(n128), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n270) );
  GTECH_FJK1S A_reg_3_ ( .J(n128), .K(n128), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n269) );
  GTECH_FJK1S A_reg_2_ ( .J(n128), .K(n128), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n268) );
  GTECH_FJK1S A_reg_1_ ( .J(n128), .K(n128), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n267) );
  GTECH_FJK1S A_reg_0_ ( .J(n128), .K(n128), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n266) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n128), .K(n128), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n128), .K(n128), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n128), .K(n128), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n128), .K(n128), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n128), .K(n128), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n128), .K(n128), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n128), .K(n128), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n128), .K(n128), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n128), .K(n128), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n128), .K(n128), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n128), .K(n128), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n128), .K(n128), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n128), .K(n128), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n128), .K(n128), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n128), .K(n128), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n128), .K(n128), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n128), .K(n128), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n128), .K(n128), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n128), .K(n128), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n128), .K(n128), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n128), .K(n128), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n128), .K(n128), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n128), .K(n128), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n128), .K(n128), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n128), .K(n128), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n128), .K(n128), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n128), .K(n128), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n128), .K(n128), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n128), .K(n128), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n128), .K(n128), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n128), .K(n128), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n128), .K(n128), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n128), .K(n128), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n128), .K(n128), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n128), .K(n128), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n128), .K(n128), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n128), .K(n128), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n128), .K(n128), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n128), .K(n128), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n128), .K(n128), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n128), .K(n128), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n128), .K(n128), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n128), .K(n128), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n128), .K(n128), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n128), .K(n128), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n128), .K(n128), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n128), .K(n128), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n128), .K(n128), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n128), .K(n128), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n128), .K(n128), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n128), .K(n128), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n128), .K(n128), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n128), .K(n128), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n128), .K(n128), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n128), .K(n128), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n128), .K(n128), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n128), .K(n128), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n128), .K(n128), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n128), .K(n128), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n128), .K(n128), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n128), .K(n128), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n128), .K(n128), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n128), .K(n128), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n128), .K(n128), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n128), .K(n128), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n128), .K(n128), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U267 ( .Z(n128) );
  GTECH_NOT U268 ( .A(n283), .Z(N99) );
  GTECH_AOI222 U269 ( .A(n284), .B(n285), .C(n286), .D(n287), .E(n288), .F(
        n289), .Z(n283) );
  GTECH_NOT U270 ( .A(n290), .Z(N98) );
  GTECH_AOI222 U271 ( .A(n286), .B(n291), .C(n292), .D(n293), .E(R[15]), .F(
        n294), .Z(n290) );
  GTECH_NAND2 U272 ( .A(n295), .B(n296), .Z(n292) );
  GTECH_AO22 U273 ( .A(n297), .B(n298), .C(R[14]), .D(n294), .Z(N97) );
  GTECH_AO22 U274 ( .A(n297), .B(n299), .C(R[13]), .D(n294), .Z(N96) );
  GTECH_AO22 U275 ( .A(n297), .B(n300), .C(R[12]), .D(n294), .Z(N95) );
  GTECH_AO22 U276 ( .A(n297), .B(n301), .C(R[11]), .D(n294), .Z(N94) );
  GTECH_AO22 U277 ( .A(n297), .B(n302), .C(R[10]), .D(n294), .Z(N93) );
  GTECH_AO22 U278 ( .A(n297), .B(n303), .C(R[9]), .D(n294), .Z(N92) );
  GTECH_AO22 U279 ( .A(n297), .B(n304), .C(R[8]), .D(n294), .Z(N91) );
  GTECH_AO22 U280 ( .A(n297), .B(n305), .C(R[7]), .D(n294), .Z(N90) );
  GTECH_AO22 U281 ( .A(n297), .B(n306), .C(R[6]), .D(n294), .Z(N89) );
  GTECH_AO22 U282 ( .A(n297), .B(n307), .C(R[5]), .D(n294), .Z(N88) );
  GTECH_AO22 U283 ( .A(n297), .B(n308), .C(R[4]), .D(n294), .Z(N87) );
  GTECH_AO22 U284 ( .A(n297), .B(n309), .C(R[3]), .D(n294), .Z(N86) );
  GTECH_AO22 U285 ( .A(n297), .B(n310), .C(R[2]), .D(n294), .Z(N85) );
  GTECH_AO22 U286 ( .A(n297), .B(n311), .C(R[1]), .D(n294), .Z(N84) );
  GTECH_AO22 U287 ( .A(n297), .B(n312), .C(R[0]), .D(n294), .Z(N83) );
  GTECH_AND2 U288 ( .A(M[15]), .B(n294), .Z(N42) );
  GTECH_AND2 U289 ( .A(M[14]), .B(n294), .Z(N39) );
  GTECH_AND2 U290 ( .A(M[13]), .B(n294), .Z(N38) );
  GTECH_AND2 U291 ( .A(M[12]), .B(n294), .Z(N37) );
  GTECH_AND2 U292 ( .A(M[11]), .B(n294), .Z(N36) );
  GTECH_AND2 U293 ( .A(M[10]), .B(n294), .Z(N35) );
  GTECH_AND2 U294 ( .A(M[9]), .B(n294), .Z(N34) );
  GTECH_AND2 U295 ( .A(M[8]), .B(n294), .Z(N33) );
  GTECH_AND2 U296 ( .A(M[7]), .B(n294), .Z(N32) );
  GTECH_AND2 U297 ( .A(M[6]), .B(n294), .Z(N31) );
  GTECH_AND2 U298 ( .A(M[5]), .B(n294), .Z(N30) );
  GTECH_AND2 U299 ( .A(M[4]), .B(n294), .Z(N29) );
  GTECH_AND2 U300 ( .A(M[3]), .B(n294), .Z(N28) );
  GTECH_AND2 U301 ( .A(M[2]), .B(n294), .Z(N27) );
  GTECH_AND2 U302 ( .A(M[1]), .B(n294), .Z(N26) );
  GTECH_AND2 U303 ( .A(M[0]), .B(n294), .Z(N25) );
  GTECH_NOT U304 ( .A(n313), .Z(n294) );
  GTECH_NAND2 U305 ( .A(n313), .B(n314), .Z(N19) );
  GTECH_NAND3 U306 ( .A(n315), .B(n316), .C(n297), .Z(n314) );
  GTECH_NAND3 U307 ( .A(n317), .B(n318), .C(n319), .Z(N18) );
  GTECH_AND2 U308 ( .A(n297), .B(n320), .Z(N17) );
  GTECH_OAI21 U309 ( .A(n8), .B(n321), .C(n315), .Z(n320) );
  GTECH_AND2 U310 ( .A(n297), .B(n322), .Z(N16) );
  GTECH_OAI21 U311 ( .A(n7), .B(n323), .C(n324), .Z(n322) );
  GTECH_NOT U312 ( .A(n325), .Z(N152) );
  GTECH_AOI222 U313 ( .A(n326), .B(n327), .C(n328), .D(n329), .E(n330), .F(
        n331), .Z(n325) );
  GTECH_NAND2 U314 ( .A(n318), .B(n332), .Z(N151) );
  GTECH_NOT U315 ( .A(n333), .Z(N150) );
  GTECH_AOI222 U316 ( .A(n334), .B(n326), .C(n328), .D(n335), .E(n330), .F(
        n336), .Z(n333) );
  GTECH_MUX2 U317 ( .A(n337), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND2 U318 ( .A(n297), .B(n338), .Z(n337) );
  GTECH_NOT U319 ( .A(n339), .Z(N149) );
  GTECH_AOI222 U320 ( .A(n340), .B(n326), .C(n328), .D(n341), .E(n330), .F(
        n342), .Z(n339) );
  GTECH_NOT U321 ( .A(n343), .Z(N148) );
  GTECH_AOI222 U322 ( .A(n344), .B(n326), .C(n328), .D(n345), .E(n330), .F(
        n346), .Z(n343) );
  GTECH_NOT U323 ( .A(n347), .Z(N147) );
  GTECH_AOI222 U324 ( .A(n348), .B(n326), .C(n328), .D(n349), .E(n330), .F(
        n350), .Z(n347) );
  GTECH_NOT U325 ( .A(n351), .Z(N146) );
  GTECH_AOI222 U326 ( .A(n352), .B(n326), .C(n328), .D(n353), .E(n330), .F(
        n354), .Z(n351) );
  GTECH_NOT U327 ( .A(n355), .Z(N145) );
  GTECH_AOI222 U328 ( .A(n356), .B(n326), .C(n328), .D(n357), .E(n330), .F(
        n358), .Z(n355) );
  GTECH_NOT U329 ( .A(n359), .Z(N144) );
  GTECH_AOI222 U330 ( .A(n360), .B(n326), .C(n328), .D(n361), .E(n330), .F(
        n362), .Z(n359) );
  GTECH_NOT U331 ( .A(n363), .Z(N143) );
  GTECH_AOI222 U332 ( .A(n364), .B(n326), .C(n328), .D(n365), .E(n330), .F(
        n366), .Z(n363) );
  GTECH_NOT U333 ( .A(n367), .Z(N142) );
  GTECH_AOI222 U334 ( .A(n368), .B(n326), .C(n328), .D(n369), .E(n330), .F(
        n370), .Z(n367) );
  GTECH_NOT U335 ( .A(n371), .Z(N141) );
  GTECH_AOI222 U336 ( .A(n372), .B(n326), .C(n328), .D(n373), .E(n330), .F(
        n374), .Z(n371) );
  GTECH_NOT U337 ( .A(n375), .Z(N140) );
  GTECH_AOI222 U338 ( .A(n376), .B(n326), .C(n328), .D(n377), .E(n330), .F(
        n378), .Z(n375) );
  GTECH_NOT U339 ( .A(n379), .Z(N14) );
  GTECH_NAND2 U340 ( .A(n297), .B(n265), .Z(n379) );
  GTECH_NOT U341 ( .A(n380), .Z(N139) );
  GTECH_AOI222 U342 ( .A(n381), .B(n326), .C(n328), .D(n382), .E(n330), .F(
        n383), .Z(n380) );
  GTECH_NOT U343 ( .A(n384), .Z(N138) );
  GTECH_AOI222 U344 ( .A(n385), .B(n326), .C(n328), .D(n386), .E(n330), .F(
        n387), .Z(n384) );
  GTECH_NOT U345 ( .A(n388), .Z(N137) );
  GTECH_AOI222 U346 ( .A(n389), .B(n326), .C(n328), .D(n390), .E(n330), .F(
        n391), .Z(n388) );
  GTECH_NOT U347 ( .A(n392), .Z(N136) );
  GTECH_AOI222 U348 ( .A(n326), .B(n285), .C(n328), .D(n287), .E(n330), .F(
        n289), .Z(n392) );
  GTECH_NOT U349 ( .A(n393), .Z(n289) );
  GTECH_XNOR2 U350 ( .A(n394), .B(n395), .Z(n393) );
  GTECH_NOT U351 ( .A(n396), .Z(n394) );
  GTECH_NOT U352 ( .A(n397), .Z(n328) );
  GTECH_NOT U353 ( .A(n398), .Z(n285) );
  GTECH_XNOR2 U354 ( .A(n399), .B(n395), .Z(n398) );
  GTECH_NOT U355 ( .A(n400), .Z(n395) );
  GTECH_XNOR2 U356 ( .A(n267), .B(n11), .Z(n400) );
  GTECH_NOT U357 ( .A(n401), .Z(n399) );
  GTECH_OAI21 U358 ( .A(n12), .B(n397), .C(n402), .Z(N135) );
  GTECH_OAI21 U359 ( .A(n330), .B(n326), .C(n293), .Z(n402) );
  GTECH_OAI21 U360 ( .A(n12), .B(n403), .C(n396), .Z(n293) );
  GTECH_NOT U361 ( .A(n404), .Z(n326) );
  GTECH_NAND3 U362 ( .A(n28), .B(n405), .C(N155), .Z(n404) );
  GTECH_NOT U363 ( .A(n406), .Z(n330) );
  GTECH_NAND3 U364 ( .A(n10), .B(n407), .C(N155), .Z(n406) );
  GTECH_NAND2 U365 ( .A(n408), .B(N155), .Z(n397) );
  GTECH_XNOR2 U366 ( .A(n28), .B(n10), .Z(n408) );
  GTECH_AND2 U367 ( .A(N155), .B(n298), .Z(N134) );
  GTECH_NOT U368 ( .A(n13), .Z(n298) );
  GTECH_AND2 U369 ( .A(N155), .B(n299), .Z(N133) );
  GTECH_NOT U370 ( .A(n14), .Z(n299) );
  GTECH_AND2 U371 ( .A(N155), .B(n300), .Z(N132) );
  GTECH_NOT U372 ( .A(n15), .Z(n300) );
  GTECH_AND2 U373 ( .A(N155), .B(n301), .Z(N131) );
  GTECH_NOT U374 ( .A(n16), .Z(n301) );
  GTECH_AND2 U375 ( .A(N155), .B(n302), .Z(N130) );
  GTECH_NOT U376 ( .A(n17), .Z(n302) );
  GTECH_AND2 U377 ( .A(N155), .B(n303), .Z(N129) );
  GTECH_NOT U378 ( .A(n18), .Z(n303) );
  GTECH_AND2 U379 ( .A(N155), .B(n304), .Z(N128) );
  GTECH_NOT U380 ( .A(n19), .Z(n304) );
  GTECH_AND2 U381 ( .A(N155), .B(n305), .Z(N127) );
  GTECH_NOT U382 ( .A(n20), .Z(n305) );
  GTECH_AND2 U383 ( .A(N155), .B(n306), .Z(N126) );
  GTECH_NOT U384 ( .A(n21), .Z(n306) );
  GTECH_AND2 U385 ( .A(N155), .B(n307), .Z(N125) );
  GTECH_NOT U386 ( .A(n22), .Z(n307) );
  GTECH_AND2 U387 ( .A(N155), .B(n308), .Z(N124) );
  GTECH_NOT U388 ( .A(n23), .Z(n308) );
  GTECH_AND2 U389 ( .A(N155), .B(n309), .Z(N123) );
  GTECH_NOT U390 ( .A(n24), .Z(n309) );
  GTECH_AND2 U391 ( .A(N155), .B(n310), .Z(N122) );
  GTECH_NOT U392 ( .A(n25), .Z(n310) );
  GTECH_AND2 U393 ( .A(N155), .B(n311), .Z(N121) );
  GTECH_NOT U394 ( .A(n26), .Z(n311) );
  GTECH_AND2 U395 ( .A(N155), .B(n312), .Z(N120) );
  GTECH_NOT U396 ( .A(n27), .Z(n312) );
  GTECH_NOT U397 ( .A(n332), .Z(N155) );
  GTECH_NAND4 U398 ( .A(n8), .B(n7), .C(n9), .D(n409), .Z(n332) );
  GTECH_AND3 U399 ( .A(n318), .B(n338), .C(n6), .Z(n409) );
  GTECH_NOT U400 ( .A(n265), .Z(n338) );
  GTECH_NOT U401 ( .A(n410), .Z(N116) );
  GTECH_AOI222 U402 ( .A(n286), .B(n329), .C(n288), .D(n331), .E(n327), .F(
        n284), .Z(n410) );
  GTECH_XNOR2 U403 ( .A(n411), .B(n412), .Z(n327) );
  GTECH_NOT U404 ( .A(n413), .Z(n412) );
  GTECH_ADD_ABC U405 ( .A(n31), .B(n281), .C(n414), .COUT(n411) );
  GTECH_XNOR2 U406 ( .A(n415), .B(n413), .Z(n331) );
  GTECH_XNOR2 U407 ( .A(n30), .B(n282), .Z(n413) );
  GTECH_AND2 U408 ( .A(n416), .B(n417), .Z(n415) );
  GTECH_OAI21 U409 ( .A(n281), .B(n335), .C(n418), .Z(n417) );
  GTECH_OR_NOT U410 ( .A(n31), .B(n281), .Z(n416) );
  GTECH_NOT U411 ( .A(n30), .Z(n329) );
  GTECH_NAND2 U412 ( .A(n319), .B(n419), .Z(N115) );
  GTECH_NOT U413 ( .A(N41), .Z(n419) );
  GTECH_NAND2 U414 ( .A(n318), .B(n313), .Z(N41) );
  GTECH_NAND2 U415 ( .A(Ld), .B(n318), .Z(n313) );
  GTECH_NOT U416 ( .A(n420), .Z(N113) );
  GTECH_AOI222 U417 ( .A(n286), .B(n335), .C(n288), .D(n336), .E(n334), .F(
        n284), .Z(n420) );
  GTECH_XNOR2 U418 ( .A(n414), .B(n421), .Z(n334) );
  GTECH_ADD_ABC U419 ( .A(n32), .B(n280), .C(n422), .COUT(n414) );
  GTECH_NOT U420 ( .A(n423), .Z(n336) );
  GTECH_XNOR2 U421 ( .A(n424), .B(n421), .Z(n423) );
  GTECH_NOT U422 ( .A(n425), .Z(n421) );
  GTECH_XNOR2 U423 ( .A(n31), .B(n281), .Z(n425) );
  GTECH_NOT U424 ( .A(n418), .Z(n424) );
  GTECH_OAI21 U425 ( .A(n32), .B(n426), .C(n427), .Z(n418) );
  GTECH_OAI21 U426 ( .A(n280), .B(n341), .C(n428), .Z(n427) );
  GTECH_NOT U427 ( .A(n280), .Z(n426) );
  GTECH_NOT U428 ( .A(n31), .Z(n335) );
  GTECH_NOT U429 ( .A(n429), .Z(N112) );
  GTECH_AOI222 U430 ( .A(n286), .B(n341), .C(n288), .D(n342), .E(n340), .F(
        n284), .Z(n429) );
  GTECH_XNOR2 U431 ( .A(n422), .B(n430), .Z(n340) );
  GTECH_ADD_ABC U432 ( .A(n33), .B(n279), .C(n431), .COUT(n422) );
  GTECH_NOT U433 ( .A(n432), .Z(n342) );
  GTECH_XNOR2 U434 ( .A(n433), .B(n430), .Z(n432) );
  GTECH_NOT U435 ( .A(n434), .Z(n430) );
  GTECH_XNOR2 U436 ( .A(n32), .B(n280), .Z(n434) );
  GTECH_NOT U437 ( .A(n428), .Z(n433) );
  GTECH_OAI21 U438 ( .A(n33), .B(n435), .C(n436), .Z(n428) );
  GTECH_OAI21 U439 ( .A(n279), .B(n345), .C(n437), .Z(n436) );
  GTECH_NOT U440 ( .A(n279), .Z(n435) );
  GTECH_NOT U441 ( .A(n32), .Z(n341) );
  GTECH_NOT U442 ( .A(n438), .Z(N111) );
  GTECH_AOI222 U443 ( .A(n286), .B(n345), .C(n288), .D(n346), .E(n344), .F(
        n284), .Z(n438) );
  GTECH_XNOR2 U444 ( .A(n431), .B(n439), .Z(n344) );
  GTECH_ADD_ABC U445 ( .A(n34), .B(n278), .C(n440), .COUT(n431) );
  GTECH_NOT U446 ( .A(n441), .Z(n346) );
  GTECH_XNOR2 U447 ( .A(n442), .B(n439), .Z(n441) );
  GTECH_NOT U448 ( .A(n443), .Z(n439) );
  GTECH_XNOR2 U449 ( .A(n33), .B(n279), .Z(n443) );
  GTECH_NOT U450 ( .A(n437), .Z(n442) );
  GTECH_OAI21 U451 ( .A(n34), .B(n444), .C(n445), .Z(n437) );
  GTECH_OAI21 U452 ( .A(n278), .B(n349), .C(n446), .Z(n445) );
  GTECH_NOT U453 ( .A(n278), .Z(n444) );
  GTECH_NOT U454 ( .A(n33), .Z(n345) );
  GTECH_NOT U455 ( .A(n447), .Z(N110) );
  GTECH_AOI222 U456 ( .A(n286), .B(n349), .C(n288), .D(n350), .E(n348), .F(
        n284), .Z(n447) );
  GTECH_XNOR2 U457 ( .A(n440), .B(n448), .Z(n348) );
  GTECH_ADD_ABC U458 ( .A(n35), .B(n277), .C(n449), .COUT(n440) );
  GTECH_NOT U459 ( .A(n450), .Z(n350) );
  GTECH_XNOR2 U460 ( .A(n451), .B(n448), .Z(n450) );
  GTECH_NOT U461 ( .A(n452), .Z(n448) );
  GTECH_XNOR2 U462 ( .A(n34), .B(n278), .Z(n452) );
  GTECH_NOT U463 ( .A(n446), .Z(n451) );
  GTECH_OAI21 U464 ( .A(n35), .B(n453), .C(n454), .Z(n446) );
  GTECH_OAI21 U465 ( .A(n277), .B(n353), .C(n455), .Z(n454) );
  GTECH_NOT U466 ( .A(n277), .Z(n453) );
  GTECH_NOT U467 ( .A(n34), .Z(n349) );
  GTECH_NOT U468 ( .A(n456), .Z(N109) );
  GTECH_AOI222 U469 ( .A(n286), .B(n353), .C(n288), .D(n354), .E(n352), .F(
        n284), .Z(n456) );
  GTECH_XNOR2 U470 ( .A(n449), .B(n457), .Z(n352) );
  GTECH_ADD_ABC U471 ( .A(n36), .B(n276), .C(n458), .COUT(n449) );
  GTECH_NOT U472 ( .A(n459), .Z(n354) );
  GTECH_XNOR2 U473 ( .A(n460), .B(n457), .Z(n459) );
  GTECH_NOT U474 ( .A(n461), .Z(n457) );
  GTECH_XNOR2 U475 ( .A(n35), .B(n277), .Z(n461) );
  GTECH_NOT U476 ( .A(n455), .Z(n460) );
  GTECH_OAI21 U477 ( .A(n36), .B(n462), .C(n463), .Z(n455) );
  GTECH_OAI21 U478 ( .A(n276), .B(n357), .C(n464), .Z(n463) );
  GTECH_NOT U479 ( .A(n276), .Z(n462) );
  GTECH_NOT U480 ( .A(n35), .Z(n353) );
  GTECH_NOT U481 ( .A(n465), .Z(N108) );
  GTECH_AOI222 U482 ( .A(n286), .B(n357), .C(n288), .D(n358), .E(n356), .F(
        n284), .Z(n465) );
  GTECH_XNOR2 U483 ( .A(n458), .B(n466), .Z(n356) );
  GTECH_ADD_ABC U484 ( .A(n37), .B(n275), .C(n467), .COUT(n458) );
  GTECH_NOT U485 ( .A(n468), .Z(n358) );
  GTECH_XNOR2 U486 ( .A(n469), .B(n466), .Z(n468) );
  GTECH_NOT U487 ( .A(n470), .Z(n466) );
  GTECH_XNOR2 U488 ( .A(n36), .B(n276), .Z(n470) );
  GTECH_NOT U489 ( .A(n464), .Z(n469) );
  GTECH_OAI21 U490 ( .A(n37), .B(n471), .C(n472), .Z(n464) );
  GTECH_OAI21 U491 ( .A(n275), .B(n361), .C(n473), .Z(n472) );
  GTECH_NOT U492 ( .A(n275), .Z(n471) );
  GTECH_NOT U493 ( .A(n36), .Z(n357) );
  GTECH_NOT U494 ( .A(n474), .Z(N107) );
  GTECH_AOI222 U495 ( .A(n286), .B(n361), .C(n288), .D(n362), .E(n360), .F(
        n284), .Z(n474) );
  GTECH_XNOR2 U496 ( .A(n467), .B(n475), .Z(n360) );
  GTECH_ADD_ABC U497 ( .A(n38), .B(n274), .C(n476), .COUT(n467) );
  GTECH_NOT U498 ( .A(n477), .Z(n362) );
  GTECH_XNOR2 U499 ( .A(n478), .B(n475), .Z(n477) );
  GTECH_NOT U500 ( .A(n479), .Z(n475) );
  GTECH_XNOR2 U501 ( .A(n37), .B(n275), .Z(n479) );
  GTECH_NOT U502 ( .A(n473), .Z(n478) );
  GTECH_OAI21 U503 ( .A(n38), .B(n480), .C(n481), .Z(n473) );
  GTECH_OAI21 U504 ( .A(n274), .B(n365), .C(n482), .Z(n481) );
  GTECH_NOT U505 ( .A(n274), .Z(n480) );
  GTECH_NOT U506 ( .A(n37), .Z(n361) );
  GTECH_NOT U507 ( .A(n483), .Z(N106) );
  GTECH_AOI222 U508 ( .A(n286), .B(n365), .C(n288), .D(n366), .E(n364), .F(
        n284), .Z(n483) );
  GTECH_XNOR2 U509 ( .A(n476), .B(n484), .Z(n364) );
  GTECH_ADD_ABC U510 ( .A(n39), .B(n273), .C(n485), .COUT(n476) );
  GTECH_NOT U511 ( .A(n486), .Z(n366) );
  GTECH_XNOR2 U512 ( .A(n487), .B(n484), .Z(n486) );
  GTECH_NOT U513 ( .A(n488), .Z(n484) );
  GTECH_XNOR2 U514 ( .A(n38), .B(n274), .Z(n488) );
  GTECH_NOT U515 ( .A(n482), .Z(n487) );
  GTECH_OAI21 U516 ( .A(n39), .B(n489), .C(n490), .Z(n482) );
  GTECH_OAI21 U517 ( .A(n273), .B(n369), .C(n491), .Z(n490) );
  GTECH_NOT U518 ( .A(n273), .Z(n489) );
  GTECH_NOT U519 ( .A(n38), .Z(n365) );
  GTECH_NOT U520 ( .A(n492), .Z(N105) );
  GTECH_AOI222 U521 ( .A(n286), .B(n369), .C(n288), .D(n370), .E(n368), .F(
        n284), .Z(n492) );
  GTECH_XNOR2 U522 ( .A(n485), .B(n493), .Z(n368) );
  GTECH_ADD_ABC U523 ( .A(n40), .B(n272), .C(n494), .COUT(n485) );
  GTECH_NOT U524 ( .A(n495), .Z(n370) );
  GTECH_XNOR2 U525 ( .A(n496), .B(n493), .Z(n495) );
  GTECH_NOT U526 ( .A(n497), .Z(n493) );
  GTECH_XNOR2 U527 ( .A(n39), .B(n273), .Z(n497) );
  GTECH_NOT U528 ( .A(n491), .Z(n496) );
  GTECH_OAI21 U529 ( .A(n40), .B(n498), .C(n499), .Z(n491) );
  GTECH_OAI21 U530 ( .A(n272), .B(n373), .C(n500), .Z(n499) );
  GTECH_NOT U531 ( .A(n272), .Z(n498) );
  GTECH_NOT U532 ( .A(n39), .Z(n369) );
  GTECH_NOT U533 ( .A(n501), .Z(N104) );
  GTECH_AOI222 U534 ( .A(n286), .B(n373), .C(n288), .D(n374), .E(n372), .F(
        n284), .Z(n501) );
  GTECH_XNOR2 U535 ( .A(n494), .B(n502), .Z(n372) );
  GTECH_ADD_ABC U536 ( .A(n41), .B(n271), .C(n503), .COUT(n494) );
  GTECH_NOT U537 ( .A(n504), .Z(n374) );
  GTECH_XNOR2 U538 ( .A(n505), .B(n502), .Z(n504) );
  GTECH_NOT U539 ( .A(n506), .Z(n502) );
  GTECH_XNOR2 U540 ( .A(n40), .B(n272), .Z(n506) );
  GTECH_NOT U541 ( .A(n500), .Z(n505) );
  GTECH_OAI21 U542 ( .A(n41), .B(n507), .C(n508), .Z(n500) );
  GTECH_OAI21 U543 ( .A(n271), .B(n377), .C(n509), .Z(n508) );
  GTECH_NOT U544 ( .A(n271), .Z(n507) );
  GTECH_NOT U545 ( .A(n40), .Z(n373) );
  GTECH_NOT U546 ( .A(n510), .Z(N103) );
  GTECH_AOI222 U547 ( .A(n286), .B(n377), .C(n288), .D(n378), .E(n376), .F(
        n284), .Z(n510) );
  GTECH_XNOR2 U548 ( .A(n503), .B(n511), .Z(n376) );
  GTECH_ADD_ABC U549 ( .A(n42), .B(n270), .C(n512), .COUT(n503) );
  GTECH_NOT U550 ( .A(n513), .Z(n378) );
  GTECH_XNOR2 U551 ( .A(n514), .B(n511), .Z(n513) );
  GTECH_NOT U552 ( .A(n515), .Z(n511) );
  GTECH_XNOR2 U553 ( .A(n41), .B(n271), .Z(n515) );
  GTECH_NOT U554 ( .A(n509), .Z(n514) );
  GTECH_OAI21 U555 ( .A(n42), .B(n516), .C(n517), .Z(n509) );
  GTECH_OAI21 U556 ( .A(n270), .B(n382), .C(n518), .Z(n517) );
  GTECH_NOT U557 ( .A(n270), .Z(n516) );
  GTECH_NOT U558 ( .A(n41), .Z(n377) );
  GTECH_NOT U559 ( .A(n519), .Z(N102) );
  GTECH_AOI222 U560 ( .A(n286), .B(n382), .C(n288), .D(n383), .E(n381), .F(
        n284), .Z(n519) );
  GTECH_XNOR2 U561 ( .A(n512), .B(n520), .Z(n381) );
  GTECH_ADD_ABC U562 ( .A(n43), .B(n269), .C(n521), .COUT(n512) );
  GTECH_NOT U563 ( .A(n522), .Z(n383) );
  GTECH_XNOR2 U564 ( .A(n523), .B(n520), .Z(n522) );
  GTECH_NOT U565 ( .A(n524), .Z(n520) );
  GTECH_XNOR2 U566 ( .A(n42), .B(n270), .Z(n524) );
  GTECH_NOT U567 ( .A(n518), .Z(n523) );
  GTECH_OAI21 U568 ( .A(n43), .B(n525), .C(n526), .Z(n518) );
  GTECH_OAI21 U569 ( .A(n269), .B(n386), .C(n527), .Z(n526) );
  GTECH_NOT U570 ( .A(n269), .Z(n525) );
  GTECH_NOT U571 ( .A(n42), .Z(n382) );
  GTECH_NOT U572 ( .A(n528), .Z(N101) );
  GTECH_AOI222 U573 ( .A(n286), .B(n386), .C(n288), .D(n387), .E(n385), .F(
        n284), .Z(n528) );
  GTECH_XNOR2 U574 ( .A(n521), .B(n529), .Z(n385) );
  GTECH_ADD_ABC U575 ( .A(n29), .B(n268), .C(n530), .COUT(n521) );
  GTECH_NOT U576 ( .A(n531), .Z(n387) );
  GTECH_XNOR2 U577 ( .A(n532), .B(n529), .Z(n531) );
  GTECH_NOT U578 ( .A(n533), .Z(n529) );
  GTECH_XNOR2 U579 ( .A(n43), .B(n269), .Z(n533) );
  GTECH_NOT U580 ( .A(n527), .Z(n532) );
  GTECH_OAI21 U581 ( .A(n29), .B(n534), .C(n535), .Z(n527) );
  GTECH_OAI21 U582 ( .A(n268), .B(n390), .C(n536), .Z(n535) );
  GTECH_NOT U583 ( .A(n268), .Z(n534) );
  GTECH_NOT U584 ( .A(n43), .Z(n386) );
  GTECH_NOT U585 ( .A(n537), .Z(N100) );
  GTECH_AOI222 U586 ( .A(n389), .B(n284), .C(n286), .D(n390), .E(n288), .F(
        n391), .Z(n537) );
  GTECH_NOT U587 ( .A(n538), .Z(n391) );
  GTECH_XNOR2 U588 ( .A(n539), .B(n540), .Z(n538) );
  GTECH_NOT U589 ( .A(n536), .Z(n539) );
  GTECH_OAI21 U590 ( .A(n11), .B(n541), .C(n542), .Z(n536) );
  GTECH_OAI21 U591 ( .A(n267), .B(n287), .C(n396), .Z(n542) );
  GTECH_NAND2 U592 ( .A(n12), .B(n403), .Z(n396) );
  GTECH_NOT U593 ( .A(n11), .Z(n287) );
  GTECH_NOT U594 ( .A(n267), .Z(n541) );
  GTECH_NOT U595 ( .A(n296), .Z(n288) );
  GTECH_NAND2 U596 ( .A(N82), .B(n10), .Z(n296) );
  GTECH_NOT U597 ( .A(n543), .Z(N82) );
  GTECH_NOT U598 ( .A(n29), .Z(n390) );
  GTECH_NOT U599 ( .A(n544), .Z(n286) );
  GTECH_MUX2 U600 ( .A(n543), .B(n545), .S(n10), .Z(n544) );
  GTECH_NAND2 U601 ( .A(n28), .B(n297), .Z(n545) );
  GTECH_NAND2 U602 ( .A(n297), .B(n407), .Z(n543) );
  GTECH_NOT U603 ( .A(n28), .Z(n407) );
  GTECH_NOT U604 ( .A(n295), .Z(n284) );
  GTECH_NAND3 U605 ( .A(n297), .B(n405), .C(n28), .Z(n295) );
  GTECH_NOT U606 ( .A(n10), .Z(n405) );
  GTECH_NOT U607 ( .A(n319), .Z(n297) );
  GTECH_OAI21 U608 ( .A(n315), .B(n316), .C(n546), .Z(n319) );
  GTECH_AND2 U609 ( .A(n317), .B(n318), .Z(n546) );
  GTECH_NOT U610 ( .A(Rst), .Z(n318) );
  GTECH_NOT U611 ( .A(Ld), .Z(n317) );
  GTECH_NOT U612 ( .A(n9), .Z(n316) );
  GTECH_NAND2 U613 ( .A(n8), .B(n321), .Z(n315) );
  GTECH_NOT U614 ( .A(n324), .Z(n321) );
  GTECH_NAND2 U615 ( .A(n7), .B(n323), .Z(n324) );
  GTECH_NOT U616 ( .A(n547), .Z(n323) );
  GTECH_NAND2 U617 ( .A(n6), .B(n265), .Z(n547) );
  GTECH_XNOR2 U618 ( .A(n530), .B(n540), .Z(n389) );
  GTECH_NOT U619 ( .A(n548), .Z(n540) );
  GTECH_XNOR2 U620 ( .A(n29), .B(n268), .Z(n548) );
  GTECH_ADD_ABC U621 ( .A(n267), .B(n11), .C(n401), .COUT(n530) );
  GTECH_NAND2 U622 ( .A(n291), .B(n403), .Z(n401) );
  GTECH_NOT U623 ( .A(n266), .Z(n403) );
  GTECH_NOT U624 ( .A(n12), .Z(n291) );
endmodule

