
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381;

  GTECH_MUX2 U134 ( .A(n273), .B(n274), .S(n275), .Z(sum[9]) );
  GTECH_XOR2 U135 ( .A(n276), .B(n277), .Z(n274) );
  GTECH_XOR2 U136 ( .A(n278), .B(n276), .Z(n273) );
  GTECH_NAND2 U137 ( .A(n279), .B(n280), .Z(n276) );
  GTECH_OAI21 U138 ( .A(n281), .B(n282), .C(n283), .Z(sum[8]) );
  GTECH_MUX2 U139 ( .A(n284), .B(n285), .S(n286), .Z(sum[7]) );
  GTECH_XNOR2 U140 ( .A(n287), .B(n288), .Z(n285) );
  GTECH_AOI21 U141 ( .A(n289), .B(n290), .C(n291), .Z(n288) );
  GTECH_XOR2 U142 ( .A(n287), .B(n292), .Z(n284) );
  GTECH_XOR2 U143 ( .A(a[7]), .B(b[7]), .Z(n287) );
  GTECH_MUX2 U144 ( .A(n293), .B(n294), .S(n286), .Z(sum[6]) );
  GTECH_XNOR2 U145 ( .A(n290), .B(n295), .Z(n294) );
  GTECH_OAI21 U146 ( .A(n296), .B(n297), .C(n298), .Z(n290) );
  GTECH_XNOR2 U147 ( .A(n295), .B(n299), .Z(n293) );
  GTECH_OR_NOT U148 ( .A(n291), .B(n289), .Z(n295) );
  GTECH_MUX2 U149 ( .A(n300), .B(n301), .S(n302), .Z(sum[5]) );
  GTECH_OR_NOT U150 ( .A(n296), .B(n298), .Z(n302) );
  GTECH_ADD_ABC U151 ( .A(n303), .B(a[4]), .C(b[4]), .COUT(n301) );
  GTECH_MUX2 U152 ( .A(n304), .B(n305), .S(n306), .Z(n303) );
  GTECH_OAI21 U153 ( .A(n307), .B(n308), .C(n309), .Z(n304) );
  GTECH_AO21 U154 ( .A(n297), .B(n286), .C(n310), .Z(n300) );
  GTECH_XOR2 U155 ( .A(n311), .B(n286), .Z(sum[4]) );
  GTECH_MUX2 U156 ( .A(n312), .B(n313), .S(n306), .Z(sum[3]) );
  GTECH_XNOR2 U157 ( .A(n314), .B(n315), .Z(n313) );
  GTECH_AOI21 U158 ( .A(n316), .B(n317), .C(n318), .Z(n315) );
  GTECH_XNOR2 U159 ( .A(n314), .B(n307), .Z(n312) );
  GTECH_XOR2 U160 ( .A(n308), .B(n319), .Z(n314) );
  GTECH_MUX2 U161 ( .A(n320), .B(n321), .S(n306), .Z(sum[2]) );
  GTECH_XNOR2 U162 ( .A(n317), .B(n322), .Z(n321) );
  GTECH_OAI21 U163 ( .A(n323), .B(n324), .C(n325), .Z(n317) );
  GTECH_XNOR2 U164 ( .A(n322), .B(n326), .Z(n320) );
  GTECH_OR_NOT U165 ( .A(n318), .B(n316), .Z(n322) );
  GTECH_MUX2 U166 ( .A(n327), .B(n328), .S(n329), .Z(sum[1]) );
  GTECH_OR_NOT U167 ( .A(n323), .B(n325), .Z(n329) );
  GTECH_OAI21 U168 ( .A(n330), .B(n306), .C(n324), .Z(n328) );
  GTECH_AO21 U169 ( .A(n306), .B(n324), .C(n330), .Z(n327) );
  GTECH_NAND2 U170 ( .A(a[0]), .B(b[0]), .Z(n324) );
  GTECH_MUX2 U171 ( .A(n331), .B(n332), .S(n333), .Z(sum[15]) );
  GTECH_XNOR2 U172 ( .A(n334), .B(n335), .Z(n332) );
  GTECH_XOR2 U173 ( .A(n334), .B(n336), .Z(n331) );
  GTECH_OA21 U174 ( .A(n337), .B(n338), .C(n339), .Z(n336) );
  GTECH_XNOR2 U175 ( .A(a[15]), .B(b[15]), .Z(n334) );
  GTECH_MUX2 U176 ( .A(n340), .B(n341), .S(n333), .Z(sum[14]) );
  GTECH_XOR2 U177 ( .A(n342), .B(n343), .Z(n341) );
  GTECH_XOR2 U178 ( .A(n337), .B(n342), .Z(n340) );
  GTECH_OR_NOT U179 ( .A(n338), .B(n339), .Z(n342) );
  GTECH_AOI21 U180 ( .A(n344), .B(n345), .C(n346), .Z(n337) );
  GTECH_MUX2 U181 ( .A(n347), .B(n348), .S(n333), .Z(sum[13]) );
  GTECH_XOR2 U182 ( .A(n349), .B(n350), .Z(n348) );
  GTECH_XNOR2 U183 ( .A(n345), .B(n349), .Z(n347) );
  GTECH_OR_NOT U184 ( .A(n346), .B(n344), .Z(n349) );
  GTECH_NAND2 U185 ( .A(n351), .B(n352), .Z(sum[12]) );
  GTECH_OAI21 U186 ( .A(n345), .B(n350), .C(n333), .Z(n352) );
  GTECH_MUX2 U187 ( .A(n353), .B(n354), .S(n275), .Z(sum[11]) );
  GTECH_XOR2 U188 ( .A(n355), .B(n356), .Z(n354) );
  GTECH_XNOR2 U189 ( .A(n355), .B(n357), .Z(n353) );
  GTECH_OA21 U190 ( .A(n358), .B(n359), .C(n360), .Z(n357) );
  GTECH_XOR2 U191 ( .A(a[11]), .B(b[11]), .Z(n355) );
  GTECH_MUX2 U192 ( .A(n361), .B(n362), .S(n275), .Z(sum[10]) );
  GTECH_NOT U193 ( .A(n282), .Z(n275) );
  GTECH_XOR2 U194 ( .A(n363), .B(n364), .Z(n362) );
  GTECH_XOR2 U195 ( .A(n359), .B(n363), .Z(n361) );
  GTECH_OR_NOT U196 ( .A(n358), .B(n360), .Z(n363) );
  GTECH_AOI21 U197 ( .A(n280), .B(n365), .C(n366), .Z(n359) );
  GTECH_NOT U198 ( .A(n367), .Z(n280) );
  GTECH_XNOR2 U199 ( .A(n306), .B(n305), .Z(sum[0]) );
  GTECH_OAI21 U200 ( .A(n368), .B(n369), .C(n351), .Z(cout) );
  GTECH_OR3 U201 ( .A(n345), .B(n350), .C(n333), .Z(n351) );
  GTECH_NOT U202 ( .A(n368), .Z(n333) );
  GTECH_AND2 U203 ( .A(b[12]), .B(a[12]), .Z(n345) );
  GTECH_AOI21 U204 ( .A(n335), .B(a[15]), .C(n370), .Z(n369) );
  GTECH_OA21 U205 ( .A(a[15]), .B(n335), .C(b[15]), .Z(n370) );
  GTECH_OAI21 U206 ( .A(n343), .B(n338), .C(n339), .Z(n335) );
  GTECH_NAND2 U207 ( .A(b[14]), .B(a[14]), .Z(n339) );
  GTECH_NOR2 U208 ( .A(b[14]), .B(a[14]), .Z(n338) );
  GTECH_AOI21 U209 ( .A(n344), .B(n371), .C(n346), .Z(n343) );
  GTECH_AND2 U210 ( .A(b[13]), .B(a[13]), .Z(n346) );
  GTECH_NOT U211 ( .A(n350), .Z(n371) );
  GTECH_NOR2 U212 ( .A(a[12]), .B(b[12]), .Z(n350) );
  GTECH_NOT U213 ( .A(n372), .Z(n344) );
  GTECH_NOR2 U214 ( .A(a[13]), .B(b[13]), .Z(n372) );
  GTECH_OA21 U215 ( .A(n282), .B(n373), .C(n283), .Z(n368) );
  GTECH_NAND2 U216 ( .A(n282), .B(n281), .Z(n283) );
  GTECH_AND2 U217 ( .A(n278), .B(n374), .Z(n281) );
  GTECH_NOT U218 ( .A(n277), .Z(n374) );
  GTECH_NOT U219 ( .A(n365), .Z(n278) );
  GTECH_AND2 U220 ( .A(b[8]), .B(a[8]), .Z(n365) );
  GTECH_OAI21 U221 ( .A(a[11]), .B(n356), .C(n375), .Z(n373) );
  GTECH_AO21 U222 ( .A(n356), .B(a[11]), .C(b[11]), .Z(n375) );
  GTECH_OAI21 U223 ( .A(n364), .B(n358), .C(n360), .Z(n356) );
  GTECH_NAND2 U224 ( .A(b[10]), .B(a[10]), .Z(n360) );
  GTECH_NOR2 U225 ( .A(b[10]), .B(a[10]), .Z(n358) );
  GTECH_OA21 U226 ( .A(n367), .B(n277), .C(n279), .Z(n364) );
  GTECH_NOT U227 ( .A(n366), .Z(n279) );
  GTECH_AND2 U228 ( .A(b[9]), .B(a[9]), .Z(n366) );
  GTECH_NOR2 U229 ( .A(a[8]), .B(b[8]), .Z(n277) );
  GTECH_NOR2 U230 ( .A(a[9]), .B(b[9]), .Z(n367) );
  GTECH_MUX2 U231 ( .A(n376), .B(n311), .S(n286), .Z(n282) );
  GTECH_MUX2 U232 ( .A(n377), .B(n378), .S(n306), .Z(n286) );
  GTECH_NOT U233 ( .A(cin), .Z(n306) );
  GTECH_NOT U234 ( .A(n305), .Z(n378) );
  GTECH_XOR2 U235 ( .A(a[0]), .B(b[0]), .Z(n305) );
  GTECH_OA21 U236 ( .A(n307), .B(n308), .C(n309), .Z(n377) );
  GTECH_AO21 U237 ( .A(n308), .B(n307), .C(n319), .Z(n309) );
  GTECH_NOT U238 ( .A(b[3]), .Z(n319) );
  GTECH_NOT U239 ( .A(a[3]), .Z(n308) );
  GTECH_AOI21 U240 ( .A(n326), .B(n316), .C(n318), .Z(n307) );
  GTECH_AND2 U241 ( .A(b[2]), .B(a[2]), .Z(n318) );
  GTECH_NOT U242 ( .A(n379), .Z(n316) );
  GTECH_NOR2 U243 ( .A(b[2]), .B(a[2]), .Z(n379) );
  GTECH_OAI21 U244 ( .A(n330), .B(n323), .C(n325), .Z(n326) );
  GTECH_NAND2 U245 ( .A(b[1]), .B(a[1]), .Z(n325) );
  GTECH_NOR2 U246 ( .A(a[1]), .B(b[1]), .Z(n323) );
  GTECH_NOR2 U247 ( .A(a[0]), .B(b[0]), .Z(n330) );
  GTECH_OR_NOT U248 ( .A(n310), .B(n297), .Z(n311) );
  GTECH_NAND2 U249 ( .A(b[4]), .B(a[4]), .Z(n297) );
  GTECH_OAI21 U250 ( .A(a[7]), .B(n292), .C(n380), .Z(n376) );
  GTECH_AO21 U251 ( .A(n292), .B(a[7]), .C(b[7]), .Z(n380) );
  GTECH_AO21 U252 ( .A(n299), .B(n289), .C(n291), .Z(n292) );
  GTECH_AND2 U253 ( .A(b[6]), .B(a[6]), .Z(n291) );
  GTECH_NOT U254 ( .A(n381), .Z(n289) );
  GTECH_NOR2 U255 ( .A(b[6]), .B(a[6]), .Z(n381) );
  GTECH_OAI21 U256 ( .A(n296), .B(n310), .C(n298), .Z(n299) );
  GTECH_NAND2 U257 ( .A(b[5]), .B(a[5]), .Z(n298) );
  GTECH_NOR2 U258 ( .A(a[4]), .B(b[4]), .Z(n310) );
  GTECH_NOR2 U259 ( .A(a[5]), .B(b[5]), .Z(n296) );
endmodule

