
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NAND2 U83 ( .A(n93), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI21 U86 ( .A(n98), .B(n99), .C(n100), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_NAND2 U88 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U89 ( .A(n104), .Z(n84) );
  GTECH_NAND2 U90 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_XOR2 U91 ( .A(n106), .B(n105), .Z(N153) );
  GTECH_NOT U92 ( .A(n107), .Z(n105) );
  GTECH_XNOR3 U93 ( .A(n108), .B(n93), .C(n109), .Z(n107) );
  GTECH_NOT U94 ( .A(n95), .Z(n109) );
  GTECH_XNOR3 U95 ( .A(n101), .B(n103), .C(n98), .Z(n95) );
  GTECH_NOT U96 ( .A(n102), .Z(n98) );
  GTECH_OAI21 U97 ( .A(n110), .B(n111), .C(n112), .Z(n102) );
  GTECH_OAI21 U98 ( .A(n113), .B(n114), .C(n115), .Z(n112) );
  GTECH_NOT U99 ( .A(n116), .Z(n103) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n116) );
  GTECH_NOT U101 ( .A(n99), .Z(n101) );
  GTECH_NAND2 U102 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U103 ( .A(n117), .B(n118), .C(n119), .COUT(n93) );
  GTECH_NOT U104 ( .A(n120), .Z(n119) );
  GTECH_XOR2 U105 ( .A(n121), .B(n122), .Z(n118) );
  GTECH_AND2 U106 ( .A(I_a[7]), .B(I_b[5]), .Z(n122) );
  GTECH_NOT U107 ( .A(n94), .Z(n108) );
  GTECH_NAND2 U108 ( .A(I_a[7]), .B(n123), .Z(n94) );
  GTECH_NOT U109 ( .A(n124), .Z(n106) );
  GTECH_NAND2 U110 ( .A(n125), .B(n126), .Z(n124) );
  GTECH_NOT U111 ( .A(n127), .Z(n126) );
  GTECH_XOR2 U112 ( .A(n127), .B(n128), .Z(N152) );
  GTECH_NOT U113 ( .A(n125), .Z(n128) );
  GTECH_XOR4 U114 ( .A(n129), .B(n121), .C(n120), .D(n117), .Z(n125) );
  GTECH_ADD_ABC U115 ( .A(n130), .B(n131), .C(n132), .COUT(n117) );
  GTECH_XNOR3 U116 ( .A(n133), .B(n134), .C(n135), .Z(n131) );
  GTECH_XNOR3 U117 ( .A(n113), .B(n115), .C(n110), .Z(n120) );
  GTECH_NOT U118 ( .A(n114), .Z(n110) );
  GTECH_OAI21 U119 ( .A(n136), .B(n137), .C(n138), .Z(n114) );
  GTECH_OAI21 U120 ( .A(n139), .B(n140), .C(n141), .Z(n138) );
  GTECH_NOT U121 ( .A(n142), .Z(n115) );
  GTECH_NAND2 U122 ( .A(I_b[7]), .B(I_a[5]), .Z(n142) );
  GTECH_NOT U123 ( .A(n111), .Z(n113) );
  GTECH_NAND2 U124 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_NOT U125 ( .A(n123), .Z(n121) );
  GTECH_OAI21 U126 ( .A(n143), .B(n144), .C(n145), .Z(n123) );
  GTECH_OAI21 U127 ( .A(n133), .B(n135), .C(n134), .Z(n145) );
  GTECH_AND2 U128 ( .A(I_a[7]), .B(I_b[5]), .Z(n129) );
  GTECH_ADD_ABC U129 ( .A(n146), .B(n147), .C(n148), .COUT(n127) );
  GTECH_OA22 U130 ( .A(n149), .B(n150), .C(n151), .D(n152), .Z(n147) );
  GTECH_OA21 U131 ( .A(n153), .B(n154), .C(n155), .Z(n146) );
  GTECH_XNOR3 U132 ( .A(n156), .B(n148), .C(n157), .Z(N151) );
  GTECH_OA21 U133 ( .A(n153), .B(n154), .C(n155), .Z(n157) );
  GTECH_OAI21 U134 ( .A(n158), .B(n159), .C(n160), .Z(n155) );
  GTECH_XOR2 U135 ( .A(n130), .B(n161), .Z(n148) );
  GTECH_XOR4 U136 ( .A(n134), .B(n143), .C(n132), .D(n133), .Z(n161) );
  GTECH_NOT U137 ( .A(n144), .Z(n133) );
  GTECH_NAND2 U138 ( .A(I_a[7]), .B(I_b[4]), .Z(n144) );
  GTECH_NOT U139 ( .A(n162), .Z(n132) );
  GTECH_XNOR3 U140 ( .A(n139), .B(n141), .C(n136), .Z(n162) );
  GTECH_NOT U141 ( .A(n140), .Z(n136) );
  GTECH_OAI21 U142 ( .A(n163), .B(n164), .C(n165), .Z(n140) );
  GTECH_OAI21 U143 ( .A(n166), .B(n167), .C(n168), .Z(n165) );
  GTECH_NOT U144 ( .A(n169), .Z(n141) );
  GTECH_NAND2 U145 ( .A(I_b[7]), .B(I_a[4]), .Z(n169) );
  GTECH_NOT U146 ( .A(n137), .Z(n139) );
  GTECH_NAND2 U147 ( .A(I_b[6]), .B(I_a[5]), .Z(n137) );
  GTECH_NOT U148 ( .A(n135), .Z(n143) );
  GTECH_OAI21 U149 ( .A(n170), .B(n171), .C(n172), .Z(n135) );
  GTECH_OAI21 U150 ( .A(n173), .B(n174), .C(n175), .Z(n172) );
  GTECH_NOT U151 ( .A(n176), .Z(n134) );
  GTECH_NAND2 U152 ( .A(I_a[6]), .B(I_b[5]), .Z(n176) );
  GTECH_ADD_ABC U153 ( .A(n177), .B(n178), .C(n179), .COUT(n130) );
  GTECH_NOT U154 ( .A(n180), .Z(n179) );
  GTECH_XNOR3 U155 ( .A(n173), .B(n175), .C(n174), .Z(n178) );
  GTECH_OA22 U156 ( .A(n149), .B(n150), .C(n151), .D(n152), .Z(n156) );
  GTECH_NOT U157 ( .A(n181), .Z(n152) );
  GTECH_NOT U158 ( .A(I_a[7]), .Z(n150) );
  GTECH_XNOR3 U159 ( .A(n153), .B(n158), .C(n160), .Z(N150) );
  GTECH_XOR2 U160 ( .A(n182), .B(n177), .Z(n160) );
  GTECH_ADD_ABC U161 ( .A(n183), .B(n184), .C(n185), .COUT(n177) );
  GTECH_NOT U162 ( .A(n186), .Z(n185) );
  GTECH_XNOR3 U163 ( .A(n187), .B(n188), .C(n189), .Z(n184) );
  GTECH_XOR4 U164 ( .A(n175), .B(n170), .C(n180), .D(n173), .Z(n182) );
  GTECH_NOT U165 ( .A(n171), .Z(n173) );
  GTECH_NAND2 U166 ( .A(I_a[6]), .B(I_b[4]), .Z(n171) );
  GTECH_XNOR3 U167 ( .A(n166), .B(n168), .C(n163), .Z(n180) );
  GTECH_NOT U168 ( .A(n167), .Z(n163) );
  GTECH_OAI21 U169 ( .A(n190), .B(n191), .C(n192), .Z(n167) );
  GTECH_OAI21 U170 ( .A(n193), .B(n194), .C(n195), .Z(n192) );
  GTECH_NOT U171 ( .A(n196), .Z(n168) );
  GTECH_NAND2 U172 ( .A(I_b[7]), .B(I_a[3]), .Z(n196) );
  GTECH_NOT U173 ( .A(n164), .Z(n166) );
  GTECH_NAND2 U174 ( .A(I_b[6]), .B(I_a[4]), .Z(n164) );
  GTECH_NOT U175 ( .A(n174), .Z(n170) );
  GTECH_OAI21 U176 ( .A(n197), .B(n198), .C(n199), .Z(n174) );
  GTECH_OAI21 U177 ( .A(n187), .B(n189), .C(n188), .Z(n199) );
  GTECH_NOT U178 ( .A(n200), .Z(n175) );
  GTECH_NAND2 U179 ( .A(I_a[5]), .B(I_b[5]), .Z(n200) );
  GTECH_NOT U180 ( .A(n154), .Z(n158) );
  GTECH_XOR2 U181 ( .A(n181), .B(n151), .Z(n154) );
  GTECH_AOI2N2 U182 ( .A(n201), .B(n202), .C(n203), .D(n204), .Z(n151) );
  GTECH_NAND2 U183 ( .A(n203), .B(n204), .Z(n202) );
  GTECH_XOR2 U184 ( .A(n205), .B(n149), .Z(n181) );
  GTECH_OA21 U185 ( .A(n206), .B(n207), .C(n208), .Z(n149) );
  GTECH_OAI21 U186 ( .A(n209), .B(n210), .C(n211), .Z(n208) );
  GTECH_NAND2 U187 ( .A(I_a[7]), .B(I_b[3]), .Z(n205) );
  GTECH_NOT U188 ( .A(n159), .Z(n153) );
  GTECH_OAI2N2 U189 ( .A(n212), .B(n213), .C(n214), .D(n215), .Z(n159) );
  GTECH_NAND2 U190 ( .A(n212), .B(n213), .Z(n215) );
  GTECH_XNOR3 U191 ( .A(n212), .B(n216), .C(n214), .Z(N149) );
  GTECH_XOR2 U192 ( .A(n217), .B(n183), .Z(n214) );
  GTECH_ADD_ABC U193 ( .A(n218), .B(n219), .C(n220), .COUT(n183) );
  GTECH_XNOR3 U194 ( .A(n221), .B(n222), .C(n223), .Z(n219) );
  GTECH_OA21 U195 ( .A(n224), .B(n225), .C(n226), .Z(n218) );
  GTECH_XOR4 U196 ( .A(n188), .B(n197), .C(n186), .D(n187), .Z(n217) );
  GTECH_NOT U197 ( .A(n198), .Z(n187) );
  GTECH_NAND2 U198 ( .A(I_a[5]), .B(I_b[4]), .Z(n198) );
  GTECH_XNOR3 U199 ( .A(n193), .B(n195), .C(n190), .Z(n186) );
  GTECH_NOT U200 ( .A(n194), .Z(n190) );
  GTECH_OAI21 U201 ( .A(n227), .B(n228), .C(n229), .Z(n194) );
  GTECH_NOT U202 ( .A(n230), .Z(n195) );
  GTECH_NAND2 U203 ( .A(I_b[7]), .B(I_a[2]), .Z(n230) );
  GTECH_NOT U204 ( .A(n191), .Z(n193) );
  GTECH_NAND2 U205 ( .A(I_b[6]), .B(I_a[3]), .Z(n191) );
  GTECH_NOT U206 ( .A(n189), .Z(n197) );
  GTECH_OAI21 U207 ( .A(n231), .B(n232), .C(n233), .Z(n189) );
  GTECH_OAI21 U208 ( .A(n221), .B(n223), .C(n222), .Z(n233) );
  GTECH_NOT U209 ( .A(n234), .Z(n188) );
  GTECH_NAND2 U210 ( .A(I_b[5]), .B(I_a[4]), .Z(n234) );
  GTECH_NOT U211 ( .A(n213), .Z(n216) );
  GTECH_XNOR3 U212 ( .A(n235), .B(n203), .C(n236), .Z(n213) );
  GTECH_NOT U213 ( .A(n201), .Z(n236) );
  GTECH_XNOR3 U214 ( .A(n209), .B(n211), .C(n206), .Z(n201) );
  GTECH_NOT U215 ( .A(n210), .Z(n206) );
  GTECH_OAI21 U216 ( .A(n237), .B(n238), .C(n239), .Z(n210) );
  GTECH_OAI21 U217 ( .A(n240), .B(n241), .C(n242), .Z(n239) );
  GTECH_NOT U218 ( .A(n243), .Z(n211) );
  GTECH_NAND2 U219 ( .A(I_a[6]), .B(I_b[3]), .Z(n243) );
  GTECH_NOT U220 ( .A(n207), .Z(n209) );
  GTECH_NAND2 U221 ( .A(I_a[7]), .B(I_b[2]), .Z(n207) );
  GTECH_ADD_ABC U222 ( .A(n244), .B(n245), .C(n246), .COUT(n203) );
  GTECH_NOT U223 ( .A(n247), .Z(n246) );
  GTECH_XOR2 U224 ( .A(n248), .B(n249), .Z(n245) );
  GTECH_AND2 U225 ( .A(I_a[7]), .B(I_b[1]), .Z(n249) );
  GTECH_NOT U226 ( .A(n204), .Z(n235) );
  GTECH_NAND2 U227 ( .A(I_a[7]), .B(n250), .Z(n204) );
  GTECH_ADD_ABC U228 ( .A(n251), .B(n252), .C(n253), .COUT(n212) );
  GTECH_XNOR3 U229 ( .A(n244), .B(n254), .C(n247), .Z(n252) );
  GTECH_XOR2 U230 ( .A(n255), .B(n251), .Z(N148) );
  GTECH_ADD_ABC U231 ( .A(n256), .B(n257), .C(n258), .COUT(n251) );
  GTECH_NOT U232 ( .A(n259), .Z(n258) );
  GTECH_XNOR3 U233 ( .A(n260), .B(n261), .C(n262), .Z(n257) );
  GTECH_XOR4 U234 ( .A(n254), .B(n244), .C(n247), .D(n253), .Z(n255) );
  GTECH_XOR2 U235 ( .A(n263), .B(n264), .Z(n253) );
  GTECH_XOR4 U236 ( .A(n222), .B(n231), .C(n220), .D(n221), .Z(n264) );
  GTECH_NOT U237 ( .A(n232), .Z(n221) );
  GTECH_NAND2 U238 ( .A(I_b[4]), .B(I_a[4]), .Z(n232) );
  GTECH_XNOR3 U239 ( .A(n265), .B(n266), .C(n267), .Z(n220) );
  GTECH_NOT U240 ( .A(n229), .Z(n267) );
  GTECH_OR3 U241 ( .A(n268), .B(n269), .C(n270), .Z(n229) );
  GTECH_NOT U242 ( .A(n228), .Z(n266) );
  GTECH_NAND2 U243 ( .A(I_b[7]), .B(I_a[1]), .Z(n228) );
  GTECH_NOT U244 ( .A(n227), .Z(n265) );
  GTECH_NAND2 U245 ( .A(I_b[6]), .B(I_a[2]), .Z(n227) );
  GTECH_NOT U246 ( .A(n223), .Z(n231) );
  GTECH_OAI21 U247 ( .A(n271), .B(n272), .C(n273), .Z(n223) );
  GTECH_OAI21 U248 ( .A(n274), .B(n275), .C(n276), .Z(n273) );
  GTECH_NOT U249 ( .A(n277), .Z(n222) );
  GTECH_NAND2 U250 ( .A(I_b[5]), .B(I_a[3]), .Z(n277) );
  GTECH_OA21 U251 ( .A(n224), .B(n225), .C(n226), .Z(n263) );
  GTECH_OAI21 U252 ( .A(n278), .B(n279), .C(n280), .Z(n226) );
  GTECH_XNOR3 U253 ( .A(n240), .B(n242), .C(n237), .Z(n247) );
  GTECH_NOT U254 ( .A(n241), .Z(n237) );
  GTECH_OAI21 U255 ( .A(n281), .B(n282), .C(n283), .Z(n241) );
  GTECH_OAI21 U256 ( .A(n284), .B(n285), .C(n286), .Z(n283) );
  GTECH_NOT U257 ( .A(n287), .Z(n242) );
  GTECH_NAND2 U258 ( .A(I_a[5]), .B(I_b[3]), .Z(n287) );
  GTECH_NOT U259 ( .A(n238), .Z(n240) );
  GTECH_NAND2 U260 ( .A(I_a[6]), .B(I_b[2]), .Z(n238) );
  GTECH_ADD_ABC U261 ( .A(n260), .B(n288), .C(n289), .COUT(n244) );
  GTECH_XNOR3 U262 ( .A(n290), .B(n291), .C(n292), .Z(n288) );
  GTECH_XOR2 U263 ( .A(n293), .B(n248), .Z(n254) );
  GTECH_NOT U264 ( .A(n250), .Z(n248) );
  GTECH_OAI21 U265 ( .A(n294), .B(n295), .C(n296), .Z(n250) );
  GTECH_OAI21 U266 ( .A(n290), .B(n292), .C(n291), .Z(n296) );
  GTECH_AND2 U267 ( .A(I_a[7]), .B(I_b[1]), .Z(n293) );
  GTECH_XOR2 U268 ( .A(n297), .B(n256), .Z(N147) );
  GTECH_ADD_ABC U269 ( .A(n298), .B(n299), .C(n300), .COUT(n256) );
  GTECH_XNOR3 U270 ( .A(n301), .B(n302), .C(n303), .Z(n299) );
  GTECH_OA21 U271 ( .A(n304), .B(n305), .C(n306), .Z(n298) );
  GTECH_XOR4 U272 ( .A(n261), .B(n289), .C(n259), .D(n260), .Z(n297) );
  GTECH_ADD_ABC U273 ( .A(n301), .B(n307), .C(n308), .COUT(n260) );
  GTECH_NOT U274 ( .A(n303), .Z(n308) );
  GTECH_XNOR3 U275 ( .A(n309), .B(n310), .C(n311), .Z(n307) );
  GTECH_XNOR3 U276 ( .A(n280), .B(n225), .C(n279), .Z(n259) );
  GTECH_NOT U277 ( .A(n224), .Z(n279) );
  GTECH_XOR2 U278 ( .A(n312), .B(n270), .Z(n224) );
  GTECH_NAND2 U279 ( .A(I_b[7]), .B(I_a[0]), .Z(n270) );
  GTECH_AND2 U280 ( .A(I_b[6]), .B(I_a[1]), .Z(n312) );
  GTECH_NOT U281 ( .A(n278), .Z(n225) );
  GTECH_XNOR3 U282 ( .A(n274), .B(n276), .C(n271), .Z(n278) );
  GTECH_NOT U283 ( .A(n275), .Z(n271) );
  GTECH_OAI21 U284 ( .A(n313), .B(n314), .C(n315), .Z(n275) );
  GTECH_NOT U285 ( .A(n316), .Z(n276) );
  GTECH_NAND2 U286 ( .A(I_b[5]), .B(I_a[2]), .Z(n316) );
  GTECH_NOT U287 ( .A(n272), .Z(n274) );
  GTECH_NAND2 U288 ( .A(I_b[4]), .B(I_a[3]), .Z(n272) );
  GTECH_NOT U289 ( .A(n317), .Z(n280) );
  GTECH_OR3 U290 ( .A(n318), .B(n319), .C(n269), .Z(n317) );
  GTECH_NOT U291 ( .A(I_b[6]), .Z(n269) );
  GTECH_NOT U292 ( .A(n262), .Z(n289) );
  GTECH_XNOR3 U293 ( .A(n284), .B(n286), .C(n281), .Z(n262) );
  GTECH_NOT U294 ( .A(n285), .Z(n281) );
  GTECH_OAI21 U295 ( .A(n320), .B(n321), .C(n322), .Z(n285) );
  GTECH_OAI21 U296 ( .A(n323), .B(n324), .C(n325), .Z(n322) );
  GTECH_NOT U297 ( .A(n326), .Z(n286) );
  GTECH_NAND2 U298 ( .A(I_b[3]), .B(I_a[4]), .Z(n326) );
  GTECH_NOT U299 ( .A(n282), .Z(n284) );
  GTECH_NAND2 U300 ( .A(I_a[5]), .B(I_b[2]), .Z(n282) );
  GTECH_NOT U301 ( .A(n327), .Z(n261) );
  GTECH_XNOR3 U302 ( .A(n290), .B(n291), .C(n294), .Z(n327) );
  GTECH_NOT U303 ( .A(n292), .Z(n294) );
  GTECH_OAI21 U304 ( .A(n328), .B(n329), .C(n330), .Z(n292) );
  GTECH_OAI21 U305 ( .A(n309), .B(n311), .C(n310), .Z(n330) );
  GTECH_NOT U306 ( .A(n331), .Z(n291) );
  GTECH_NAND2 U307 ( .A(I_a[6]), .B(I_b[1]), .Z(n331) );
  GTECH_NOT U308 ( .A(n295), .Z(n290) );
  GTECH_NAND2 U309 ( .A(I_a[7]), .B(I_b[0]), .Z(n295) );
  GTECH_XOR2 U310 ( .A(n332), .B(n333), .Z(N146) );
  GTECH_OA21 U311 ( .A(n304), .B(n305), .C(n306), .Z(n333) );
  GTECH_OAI21 U312 ( .A(n334), .B(n335), .C(n336), .Z(n306) );
  GTECH_XOR4 U313 ( .A(n302), .B(n301), .C(n303), .D(n300), .Z(n332) );
  GTECH_XOR2 U314 ( .A(n318), .B(n337), .Z(n300) );
  GTECH_AND2 U315 ( .A(I_b[6]), .B(I_a[0]), .Z(n337) );
  GTECH_XNOR3 U316 ( .A(n338), .B(n339), .C(n340), .Z(n318) );
  GTECH_NOT U317 ( .A(n315), .Z(n340) );
  GTECH_OR3 U318 ( .A(n268), .B(n341), .C(n342), .Z(n315) );
  GTECH_NOT U319 ( .A(n314), .Z(n339) );
  GTECH_NAND2 U320 ( .A(I_b[5]), .B(I_a[1]), .Z(n314) );
  GTECH_NOT U321 ( .A(n313), .Z(n338) );
  GTECH_NAND2 U322 ( .A(I_b[4]), .B(I_a[2]), .Z(n313) );
  GTECH_XNOR3 U323 ( .A(n323), .B(n325), .C(n320), .Z(n303) );
  GTECH_NOT U324 ( .A(n324), .Z(n320) );
  GTECH_OAI21 U325 ( .A(n343), .B(n344), .C(n345), .Z(n324) );
  GTECH_OAI21 U326 ( .A(n346), .B(n347), .C(n348), .Z(n345) );
  GTECH_NOT U327 ( .A(n349), .Z(n325) );
  GTECH_NAND2 U328 ( .A(I_b[3]), .B(I_a[3]), .Z(n349) );
  GTECH_NOT U329 ( .A(n321), .Z(n323) );
  GTECH_NAND2 U330 ( .A(I_b[2]), .B(I_a[4]), .Z(n321) );
  GTECH_ADD_ABC U331 ( .A(n350), .B(n351), .C(n352), .COUT(n301) );
  GTECH_NOT U332 ( .A(n353), .Z(n352) );
  GTECH_XNOR3 U333 ( .A(n354), .B(n355), .C(n356), .Z(n351) );
  GTECH_NOT U334 ( .A(n357), .Z(n302) );
  GTECH_XNOR3 U335 ( .A(n309), .B(n310), .C(n328), .Z(n357) );
  GTECH_NOT U336 ( .A(n311), .Z(n328) );
  GTECH_OAI21 U337 ( .A(n358), .B(n359), .C(n360), .Z(n311) );
  GTECH_OAI21 U338 ( .A(n354), .B(n356), .C(n355), .Z(n360) );
  GTECH_NOT U339 ( .A(n361), .Z(n310) );
  GTECH_NAND2 U340 ( .A(I_a[5]), .B(I_b[1]), .Z(n361) );
  GTECH_NOT U341 ( .A(n329), .Z(n309) );
  GTECH_NAND2 U342 ( .A(I_a[6]), .B(I_b[0]), .Z(n329) );
  GTECH_XNOR3 U343 ( .A(n336), .B(n305), .C(n335), .Z(N145) );
  GTECH_NOT U344 ( .A(n304), .Z(n335) );
  GTECH_XOR2 U345 ( .A(n362), .B(n342), .Z(n304) );
  GTECH_NAND2 U346 ( .A(I_b[5]), .B(I_a[0]), .Z(n342) );
  GTECH_AND2 U347 ( .A(I_b[4]), .B(I_a[1]), .Z(n362) );
  GTECH_NOT U348 ( .A(n334), .Z(n305) );
  GTECH_XOR2 U349 ( .A(n363), .B(n350), .Z(n334) );
  GTECH_ADD_ABC U350 ( .A(n364), .B(n365), .C(n366), .COUT(n350) );
  GTECH_XNOR3 U351 ( .A(n367), .B(n368), .C(n369), .Z(n365) );
  GTECH_OA21 U352 ( .A(n370), .B(n371), .C(n372), .Z(n364) );
  GTECH_XOR4 U353 ( .A(n355), .B(n358), .C(n353), .D(n354), .Z(n363) );
  GTECH_NOT U354 ( .A(n359), .Z(n354) );
  GTECH_NAND2 U355 ( .A(I_a[5]), .B(I_b[0]), .Z(n359) );
  GTECH_XNOR3 U356 ( .A(n346), .B(n348), .C(n343), .Z(n353) );
  GTECH_NOT U357 ( .A(n347), .Z(n343) );
  GTECH_OAI21 U358 ( .A(n373), .B(n374), .C(n375), .Z(n347) );
  GTECH_NOT U359 ( .A(n376), .Z(n348) );
  GTECH_NAND2 U360 ( .A(I_b[3]), .B(I_a[2]), .Z(n376) );
  GTECH_NOT U361 ( .A(n344), .Z(n346) );
  GTECH_NAND2 U362 ( .A(I_b[2]), .B(I_a[3]), .Z(n344) );
  GTECH_NOT U363 ( .A(n356), .Z(n358) );
  GTECH_OAI21 U364 ( .A(n377), .B(n378), .C(n379), .Z(n356) );
  GTECH_OAI21 U365 ( .A(n367), .B(n369), .C(n368), .Z(n379) );
  GTECH_NOT U366 ( .A(n380), .Z(n355) );
  GTECH_NAND2 U367 ( .A(I_a[4]), .B(I_b[1]), .Z(n380) );
  GTECH_NOT U368 ( .A(n381), .Z(n336) );
  GTECH_OR3 U369 ( .A(n382), .B(n319), .C(n341), .Z(n381) );
  GTECH_NOT U370 ( .A(I_b[4]), .Z(n341) );
  GTECH_XOR2 U371 ( .A(n383), .B(n382), .Z(N144) );
  GTECH_XOR2 U372 ( .A(n384), .B(n385), .Z(n382) );
  GTECH_XOR4 U373 ( .A(n368), .B(n377), .C(n366), .D(n367), .Z(n385) );
  GTECH_NOT U374 ( .A(n378), .Z(n367) );
  GTECH_NAND2 U375 ( .A(I_a[4]), .B(I_b[0]), .Z(n378) );
  GTECH_XNOR3 U376 ( .A(n386), .B(n387), .C(n388), .Z(n366) );
  GTECH_NOT U377 ( .A(n375), .Z(n388) );
  GTECH_OR3 U378 ( .A(n268), .B(n389), .C(n390), .Z(n375) );
  GTECH_NOT U379 ( .A(n374), .Z(n387) );
  GTECH_NAND2 U380 ( .A(I_b[3]), .B(I_a[1]), .Z(n374) );
  GTECH_NOT U381 ( .A(n373), .Z(n386) );
  GTECH_NAND2 U382 ( .A(I_b[2]), .B(I_a[2]), .Z(n373) );
  GTECH_NOT U383 ( .A(n369), .Z(n377) );
  GTECH_OAI21 U384 ( .A(n391), .B(n392), .C(n393), .Z(n369) );
  GTECH_OAI21 U385 ( .A(n394), .B(n395), .C(n396), .Z(n393) );
  GTECH_NOT U386 ( .A(n397), .Z(n368) );
  GTECH_NAND2 U387 ( .A(I_a[3]), .B(I_b[1]), .Z(n397) );
  GTECH_OA21 U388 ( .A(n370), .B(n371), .C(n372), .Z(n384) );
  GTECH_OAI21 U389 ( .A(n398), .B(n399), .C(n400), .Z(n372) );
  GTECH_NAND2 U390 ( .A(I_b[4]), .B(I_a[0]), .Z(n383) );
  GTECH_XNOR3 U391 ( .A(n400), .B(n371), .C(n399), .Z(N143) );
  GTECH_NOT U392 ( .A(n370), .Z(n399) );
  GTECH_XOR2 U393 ( .A(n401), .B(n390), .Z(n370) );
  GTECH_NAND2 U394 ( .A(I_b[3]), .B(I_a[0]), .Z(n390) );
  GTECH_AND2 U395 ( .A(I_b[2]), .B(I_a[1]), .Z(n401) );
  GTECH_NOT U396 ( .A(n398), .Z(n371) );
  GTECH_XNOR3 U397 ( .A(n394), .B(n396), .C(n391), .Z(n398) );
  GTECH_NOT U398 ( .A(n395), .Z(n391) );
  GTECH_OAI21 U399 ( .A(n402), .B(n403), .C(n404), .Z(n395) );
  GTECH_NOT U400 ( .A(n405), .Z(n396) );
  GTECH_NAND2 U401 ( .A(I_b[1]), .B(I_a[2]), .Z(n405) );
  GTECH_NOT U402 ( .A(n392), .Z(n394) );
  GTECH_NAND2 U403 ( .A(I_b[0]), .B(I_a[3]), .Z(n392) );
  GTECH_NOT U404 ( .A(n406), .Z(n400) );
  GTECH_OR3 U405 ( .A(n407), .B(n319), .C(n389), .Z(n406) );
  GTECH_NOT U406 ( .A(I_b[2]), .Z(n389) );
  GTECH_NOT U407 ( .A(I_a[0]), .Z(n319) );
  GTECH_XOR2 U408 ( .A(n408), .B(n407), .Z(N142) );
  GTECH_XNOR3 U409 ( .A(n409), .B(n410), .C(n411), .Z(n407) );
  GTECH_NOT U410 ( .A(n404), .Z(n411) );
  GTECH_OR3 U411 ( .A(n412), .B(n413), .C(n268), .Z(n404) );
  GTECH_NOT U412 ( .A(I_a[1]), .Z(n268) );
  GTECH_NOT U413 ( .A(I_b[0]), .Z(n412) );
  GTECH_NOT U414 ( .A(n402), .Z(n410) );
  GTECH_NAND2 U415 ( .A(I_a[1]), .B(I_b[1]), .Z(n402) );
  GTECH_NOT U416 ( .A(n403), .Z(n409) );
  GTECH_NAND2 U417 ( .A(I_b[0]), .B(I_a[2]), .Z(n403) );
  GTECH_NAND2 U418 ( .A(I_b[2]), .B(I_a[0]), .Z(n408) );
  GTECH_XOR2 U419 ( .A(n414), .B(n413), .Z(N141) );
  GTECH_NAND2 U420 ( .A(I_a[0]), .B(I_b[1]), .Z(n413) );
  GTECH_NAND2 U421 ( .A(I_a[1]), .B(I_b[0]), .Z(n414) );
  GTECH_AND2 U422 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

