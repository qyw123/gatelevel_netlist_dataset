
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NAND2 U83 ( .A(n93), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI21 U86 ( .A(n98), .B(n99), .C(n100), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_NAND2 U88 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U89 ( .A(n104), .Z(n84) );
  GTECH_NAND2 U90 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_XOR2 U91 ( .A(n106), .B(n105), .Z(N153) );
  GTECH_NOT U92 ( .A(n107), .Z(n105) );
  GTECH_XNOR3 U93 ( .A(n108), .B(n93), .C(n109), .Z(n107) );
  GTECH_NOT U94 ( .A(n95), .Z(n109) );
  GTECH_XNOR3 U95 ( .A(n101), .B(n103), .C(n98), .Z(n95) );
  GTECH_NOT U96 ( .A(n102), .Z(n98) );
  GTECH_OAI21 U97 ( .A(n110), .B(n111), .C(n112), .Z(n102) );
  GTECH_OAI21 U98 ( .A(n113), .B(n114), .C(n115), .Z(n112) );
  GTECH_NOT U99 ( .A(n116), .Z(n103) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n116) );
  GTECH_NOT U101 ( .A(n99), .Z(n101) );
  GTECH_NAND2 U102 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U103 ( .A(n117), .B(n118), .C(n119), .COUT(n93) );
  GTECH_XOR2 U104 ( .A(n120), .B(n121), .Z(n118) );
  GTECH_AND2 U105 ( .A(I_a[7]), .B(I_b[5]), .Z(n121) );
  GTECH_NOT U106 ( .A(n94), .Z(n108) );
  GTECH_NAND2 U107 ( .A(I_a[7]), .B(n122), .Z(n94) );
  GTECH_NOT U108 ( .A(n123), .Z(n106) );
  GTECH_NAND2 U109 ( .A(n124), .B(n125), .Z(n123) );
  GTECH_NOT U110 ( .A(n126), .Z(n125) );
  GTECH_XOR2 U111 ( .A(n126), .B(n127), .Z(N152) );
  GTECH_NOT U112 ( .A(n124), .Z(n127) );
  GTECH_XNOR4 U113 ( .A(n128), .B(n120), .C(n117), .D(n119), .Z(n124) );
  GTECH_NOT U114 ( .A(n129), .Z(n119) );
  GTECH_XNOR3 U115 ( .A(n113), .B(n115), .C(n110), .Z(n129) );
  GTECH_NOT U116 ( .A(n114), .Z(n110) );
  GTECH_OAI21 U117 ( .A(n130), .B(n131), .C(n132), .Z(n114) );
  GTECH_OAI21 U118 ( .A(n133), .B(n134), .C(n135), .Z(n132) );
  GTECH_NOT U119 ( .A(n136), .Z(n115) );
  GTECH_NAND2 U120 ( .A(I_b[7]), .B(I_a[5]), .Z(n136) );
  GTECH_NOT U121 ( .A(n111), .Z(n113) );
  GTECH_NAND2 U122 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_ADD_ABC U123 ( .A(n137), .B(n138), .C(n139), .COUT(n117) );
  GTECH_NOT U124 ( .A(n140), .Z(n139) );
  GTECH_XNOR3 U125 ( .A(n141), .B(n142), .C(n143), .Z(n138) );
  GTECH_NOT U126 ( .A(n122), .Z(n120) );
  GTECH_OAI21 U127 ( .A(n144), .B(n145), .C(n146), .Z(n122) );
  GTECH_OAI21 U128 ( .A(n141), .B(n143), .C(n142), .Z(n146) );
  GTECH_AND2 U129 ( .A(I_a[7]), .B(I_b[5]), .Z(n128) );
  GTECH_ADD_ABC U130 ( .A(n147), .B(n148), .C(n149), .COUT(n126) );
  GTECH_OA22 U131 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n148) );
  GTECH_OA21 U132 ( .A(n154), .B(n155), .C(n156), .Z(n147) );
  GTECH_XNOR3 U133 ( .A(n157), .B(n149), .C(n158), .Z(N151) );
  GTECH_OA21 U134 ( .A(n154), .B(n155), .C(n156), .Z(n158) );
  GTECH_OAI21 U135 ( .A(n159), .B(n160), .C(n161), .Z(n156) );
  GTECH_XOR2 U136 ( .A(n137), .B(n162), .Z(n149) );
  GTECH_XNOR4 U137 ( .A(n142), .B(n144), .C(n140), .D(n141), .Z(n162) );
  GTECH_NOT U138 ( .A(n145), .Z(n141) );
  GTECH_NAND2 U139 ( .A(I_a[7]), .B(I_b[4]), .Z(n145) );
  GTECH_XNOR3 U140 ( .A(n133), .B(n135), .C(n130), .Z(n140) );
  GTECH_NOT U141 ( .A(n134), .Z(n130) );
  GTECH_OAI21 U142 ( .A(n163), .B(n164), .C(n165), .Z(n134) );
  GTECH_OAI21 U143 ( .A(n166), .B(n167), .C(n168), .Z(n165) );
  GTECH_NOT U144 ( .A(n169), .Z(n135) );
  GTECH_NAND2 U145 ( .A(I_b[7]), .B(I_a[4]), .Z(n169) );
  GTECH_NOT U146 ( .A(n131), .Z(n133) );
  GTECH_NAND2 U147 ( .A(I_b[6]), .B(I_a[5]), .Z(n131) );
  GTECH_NOT U148 ( .A(n143), .Z(n144) );
  GTECH_OAI21 U149 ( .A(n170), .B(n171), .C(n172), .Z(n143) );
  GTECH_OAI21 U150 ( .A(n173), .B(n174), .C(n175), .Z(n172) );
  GTECH_NOT U151 ( .A(n176), .Z(n142) );
  GTECH_NAND2 U152 ( .A(I_a[6]), .B(I_b[5]), .Z(n176) );
  GTECH_ADD_ABC U153 ( .A(n177), .B(n178), .C(n179), .COUT(n137) );
  GTECH_XNOR3 U154 ( .A(n173), .B(n175), .C(n174), .Z(n178) );
  GTECH_OA22 U155 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n157) );
  GTECH_NOT U156 ( .A(n180), .Z(n153) );
  GTECH_NOT U157 ( .A(I_a[7]), .Z(n151) );
  GTECH_XNOR3 U158 ( .A(n154), .B(n159), .C(n161), .Z(N150) );
  GTECH_XOR2 U159 ( .A(n181), .B(n177), .Z(n161) );
  GTECH_ADD_ABC U160 ( .A(n182), .B(n183), .C(n184), .COUT(n177) );
  GTECH_XNOR3 U161 ( .A(n185), .B(n186), .C(n187), .Z(n183) );
  GTECH_XNOR4 U162 ( .A(n175), .B(n170), .C(n179), .D(n173), .Z(n181) );
  GTECH_NOT U163 ( .A(n171), .Z(n173) );
  GTECH_NAND2 U164 ( .A(I_a[6]), .B(I_b[4]), .Z(n171) );
  GTECH_NOT U165 ( .A(n188), .Z(n179) );
  GTECH_XNOR3 U166 ( .A(n166), .B(n168), .C(n163), .Z(n188) );
  GTECH_NOT U167 ( .A(n167), .Z(n163) );
  GTECH_OAI21 U168 ( .A(n189), .B(n190), .C(n191), .Z(n167) );
  GTECH_OAI21 U169 ( .A(n192), .B(n193), .C(n194), .Z(n191) );
  GTECH_NOT U170 ( .A(n195), .Z(n168) );
  GTECH_NAND2 U171 ( .A(I_b[7]), .B(I_a[3]), .Z(n195) );
  GTECH_NOT U172 ( .A(n164), .Z(n166) );
  GTECH_NAND2 U173 ( .A(I_b[6]), .B(I_a[4]), .Z(n164) );
  GTECH_NOT U174 ( .A(n174), .Z(n170) );
  GTECH_OAI21 U175 ( .A(n196), .B(n197), .C(n198), .Z(n174) );
  GTECH_OAI21 U176 ( .A(n185), .B(n187), .C(n186), .Z(n198) );
  GTECH_NOT U177 ( .A(n199), .Z(n175) );
  GTECH_NAND2 U178 ( .A(I_a[5]), .B(I_b[5]), .Z(n199) );
  GTECH_NOT U179 ( .A(n155), .Z(n159) );
  GTECH_XOR2 U180 ( .A(n180), .B(n152), .Z(n155) );
  GTECH_AOI2N2 U181 ( .A(n200), .B(n201), .C(n202), .D(n203), .Z(n152) );
  GTECH_NAND2 U182 ( .A(n202), .B(n203), .Z(n201) );
  GTECH_XOR2 U183 ( .A(n204), .B(n150), .Z(n180) );
  GTECH_OA21 U184 ( .A(n205), .B(n206), .C(n207), .Z(n150) );
  GTECH_OAI21 U185 ( .A(n208), .B(n209), .C(n210), .Z(n207) );
  GTECH_NAND2 U186 ( .A(I_a[7]), .B(I_b[3]), .Z(n204) );
  GTECH_NOT U187 ( .A(n160), .Z(n154) );
  GTECH_OAI2N2 U188 ( .A(n211), .B(n212), .C(n213), .D(n214), .Z(n160) );
  GTECH_NAND2 U189 ( .A(n211), .B(n212), .Z(n214) );
  GTECH_XNOR3 U190 ( .A(n211), .B(n215), .C(n213), .Z(N149) );
  GTECH_XOR2 U191 ( .A(n216), .B(n182), .Z(n213) );
  GTECH_ADD_ABC U192 ( .A(n217), .B(n218), .C(n219), .COUT(n182) );
  GTECH_XNOR3 U193 ( .A(n220), .B(n221), .C(n222), .Z(n218) );
  GTECH_OA21 U194 ( .A(n223), .B(n224), .C(n225), .Z(n217) );
  GTECH_XNOR4 U195 ( .A(n186), .B(n196), .C(n184), .D(n185), .Z(n216) );
  GTECH_NOT U196 ( .A(n197), .Z(n185) );
  GTECH_NAND2 U197 ( .A(I_a[5]), .B(I_b[4]), .Z(n197) );
  GTECH_NOT U198 ( .A(n226), .Z(n184) );
  GTECH_XNOR3 U199 ( .A(n192), .B(n194), .C(n189), .Z(n226) );
  GTECH_NOT U200 ( .A(n193), .Z(n189) );
  GTECH_OAI21 U201 ( .A(n227), .B(n228), .C(n229), .Z(n193) );
  GTECH_NOT U202 ( .A(n230), .Z(n194) );
  GTECH_NAND2 U203 ( .A(I_b[7]), .B(I_a[2]), .Z(n230) );
  GTECH_NOT U204 ( .A(n190), .Z(n192) );
  GTECH_NAND2 U205 ( .A(I_b[6]), .B(I_a[3]), .Z(n190) );
  GTECH_NOT U206 ( .A(n187), .Z(n196) );
  GTECH_OAI21 U207 ( .A(n231), .B(n232), .C(n233), .Z(n187) );
  GTECH_OAI21 U208 ( .A(n220), .B(n222), .C(n221), .Z(n233) );
  GTECH_NOT U209 ( .A(n232), .Z(n220) );
  GTECH_NOT U210 ( .A(n234), .Z(n186) );
  GTECH_NAND2 U211 ( .A(I_b[5]), .B(I_a[4]), .Z(n234) );
  GTECH_NOT U212 ( .A(n212), .Z(n215) );
  GTECH_XNOR3 U213 ( .A(n235), .B(n202), .C(n236), .Z(n212) );
  GTECH_NOT U214 ( .A(n200), .Z(n236) );
  GTECH_XNOR3 U215 ( .A(n208), .B(n210), .C(n205), .Z(n200) );
  GTECH_NOT U216 ( .A(n209), .Z(n205) );
  GTECH_OAI21 U217 ( .A(n237), .B(n238), .C(n239), .Z(n209) );
  GTECH_OAI21 U218 ( .A(n240), .B(n241), .C(n242), .Z(n239) );
  GTECH_NOT U219 ( .A(n243), .Z(n210) );
  GTECH_NAND2 U220 ( .A(I_a[6]), .B(I_b[3]), .Z(n243) );
  GTECH_NOT U221 ( .A(n206), .Z(n208) );
  GTECH_NAND2 U222 ( .A(I_a[7]), .B(I_b[2]), .Z(n206) );
  GTECH_ADD_ABC U223 ( .A(n244), .B(n245), .C(n246), .COUT(n202) );
  GTECH_XOR2 U224 ( .A(n247), .B(n248), .Z(n245) );
  GTECH_AND2 U225 ( .A(I_a[7]), .B(I_b[1]), .Z(n248) );
  GTECH_NOT U226 ( .A(n203), .Z(n235) );
  GTECH_NAND2 U227 ( .A(I_a[7]), .B(n249), .Z(n203) );
  GTECH_ADD_ABC U228 ( .A(n250), .B(n251), .C(n252), .COUT(n211) );
  GTECH_XNOR3 U229 ( .A(n244), .B(n253), .C(n254), .Z(n251) );
  GTECH_XOR2 U230 ( .A(n255), .B(n250), .Z(N148) );
  GTECH_ADD_ABC U231 ( .A(n256), .B(n257), .C(n258), .COUT(n250) );
  GTECH_XNOR3 U232 ( .A(n259), .B(n260), .C(n261), .Z(n257) );
  GTECH_XNOR4 U233 ( .A(n253), .B(n246), .C(n252), .D(n244), .Z(n255) );
  GTECH_ADD_ABC U234 ( .A(n259), .B(n262), .C(n263), .COUT(n244) );
  GTECH_XNOR3 U235 ( .A(n264), .B(n265), .C(n266), .Z(n262) );
  GTECH_XOR2 U236 ( .A(n267), .B(n268), .Z(n252) );
  GTECH_XNOR4 U237 ( .A(n221), .B(n231), .C(n232), .D(n219), .Z(n268) );
  GTECH_XNOR3 U238 ( .A(n269), .B(n270), .C(n271), .Z(n219) );
  GTECH_NOT U239 ( .A(n229), .Z(n271) );
  GTECH_NAND3 U240 ( .A(I_b[6]), .B(I_a[1]), .C(n272), .Z(n229) );
  GTECH_NOT U241 ( .A(n228), .Z(n270) );
  GTECH_NAND2 U242 ( .A(I_b[7]), .B(I_a[1]), .Z(n228) );
  GTECH_NOT U243 ( .A(n227), .Z(n269) );
  GTECH_NAND2 U244 ( .A(I_b[6]), .B(I_a[2]), .Z(n227) );
  GTECH_NAND2 U245 ( .A(I_b[4]), .B(I_a[4]), .Z(n232) );
  GTECH_NOT U246 ( .A(n222), .Z(n231) );
  GTECH_OAI21 U247 ( .A(n273), .B(n274), .C(n275), .Z(n222) );
  GTECH_OAI21 U248 ( .A(n276), .B(n277), .C(n278), .Z(n275) );
  GTECH_NOT U249 ( .A(n279), .Z(n221) );
  GTECH_NAND2 U250 ( .A(I_b[5]), .B(I_a[3]), .Z(n279) );
  GTECH_OA21 U251 ( .A(n223), .B(n224), .C(n225), .Z(n267) );
  GTECH_OAI21 U252 ( .A(n280), .B(n281), .C(n282), .Z(n225) );
  GTECH_NOT U253 ( .A(n254), .Z(n246) );
  GTECH_XNOR3 U254 ( .A(n240), .B(n242), .C(n237), .Z(n254) );
  GTECH_NOT U255 ( .A(n241), .Z(n237) );
  GTECH_OAI21 U256 ( .A(n283), .B(n284), .C(n285), .Z(n241) );
  GTECH_OAI21 U257 ( .A(n286), .B(n287), .C(n288), .Z(n285) );
  GTECH_NOT U258 ( .A(n289), .Z(n242) );
  GTECH_NAND2 U259 ( .A(I_a[5]), .B(I_b[3]), .Z(n289) );
  GTECH_NOT U260 ( .A(n238), .Z(n240) );
  GTECH_NAND2 U261 ( .A(I_a[6]), .B(I_b[2]), .Z(n238) );
  GTECH_XOR2 U262 ( .A(n290), .B(n247), .Z(n253) );
  GTECH_NOT U263 ( .A(n249), .Z(n247) );
  GTECH_OAI21 U264 ( .A(n291), .B(n292), .C(n293), .Z(n249) );
  GTECH_OAI21 U265 ( .A(n264), .B(n266), .C(n265), .Z(n293) );
  GTECH_AND2 U266 ( .A(I_a[7]), .B(I_b[1]), .Z(n290) );
  GTECH_XOR2 U267 ( .A(n294), .B(n256), .Z(N147) );
  GTECH_ADD_ABC U268 ( .A(n295), .B(n296), .C(n297), .COUT(n256) );
  GTECH_XNOR3 U269 ( .A(n298), .B(n299), .C(n300), .Z(n296) );
  GTECH_OA21 U270 ( .A(n301), .B(n302), .C(n303), .Z(n295) );
  GTECH_XNOR4 U271 ( .A(n260), .B(n263), .C(n258), .D(n259), .Z(n294) );
  GTECH_ADD_ABC U272 ( .A(n298), .B(n304), .C(n305), .COUT(n259) );
  GTECH_XNOR3 U273 ( .A(n306), .B(n307), .C(n308), .Z(n304) );
  GTECH_NOT U274 ( .A(n309), .Z(n258) );
  GTECH_XNOR3 U275 ( .A(n282), .B(n224), .C(n281), .Z(n309) );
  GTECH_NOT U276 ( .A(n223), .Z(n281) );
  GTECH_XOR2 U277 ( .A(n310), .B(n272), .Z(n223) );
  GTECH_NOT U278 ( .A(n311), .Z(n272) );
  GTECH_NAND2 U279 ( .A(I_b[7]), .B(I_a[0]), .Z(n311) );
  GTECH_NAND2 U280 ( .A(I_b[6]), .B(I_a[1]), .Z(n310) );
  GTECH_NOT U281 ( .A(n280), .Z(n224) );
  GTECH_XNOR3 U282 ( .A(n276), .B(n278), .C(n273), .Z(n280) );
  GTECH_NOT U283 ( .A(n277), .Z(n273) );
  GTECH_OAI21 U284 ( .A(n312), .B(n313), .C(n314), .Z(n277) );
  GTECH_NOT U285 ( .A(n315), .Z(n278) );
  GTECH_NAND2 U286 ( .A(I_b[5]), .B(I_a[2]), .Z(n315) );
  GTECH_NOT U287 ( .A(n274), .Z(n276) );
  GTECH_NAND2 U288 ( .A(I_b[4]), .B(I_a[3]), .Z(n274) );
  GTECH_NOT U289 ( .A(n316), .Z(n282) );
  GTECH_NAND3 U290 ( .A(I_a[0]), .B(n317), .C(I_b[6]), .Z(n316) );
  GTECH_NOT U291 ( .A(n318), .Z(n317) );
  GTECH_NOT U292 ( .A(n261), .Z(n263) );
  GTECH_XNOR3 U293 ( .A(n286), .B(n288), .C(n283), .Z(n261) );
  GTECH_NOT U294 ( .A(n287), .Z(n283) );
  GTECH_OAI21 U295 ( .A(n319), .B(n320), .C(n321), .Z(n287) );
  GTECH_OAI21 U296 ( .A(n322), .B(n323), .C(n324), .Z(n321) );
  GTECH_NOT U297 ( .A(n325), .Z(n288) );
  GTECH_NAND2 U298 ( .A(I_b[3]), .B(I_a[4]), .Z(n325) );
  GTECH_NOT U299 ( .A(n284), .Z(n286) );
  GTECH_NAND2 U300 ( .A(I_a[5]), .B(I_b[2]), .Z(n284) );
  GTECH_NOT U301 ( .A(n326), .Z(n260) );
  GTECH_XNOR3 U302 ( .A(n264), .B(n265), .C(n291), .Z(n326) );
  GTECH_NOT U303 ( .A(n266), .Z(n291) );
  GTECH_OAI21 U304 ( .A(n327), .B(n328), .C(n329), .Z(n266) );
  GTECH_OAI21 U305 ( .A(n306), .B(n308), .C(n307), .Z(n329) );
  GTECH_NOT U306 ( .A(n330), .Z(n265) );
  GTECH_NAND2 U307 ( .A(I_a[6]), .B(I_b[1]), .Z(n330) );
  GTECH_NOT U308 ( .A(n292), .Z(n264) );
  GTECH_NAND2 U309 ( .A(I_a[7]), .B(I_b[0]), .Z(n292) );
  GTECH_XOR2 U310 ( .A(n331), .B(n332), .Z(N146) );
  GTECH_OA21 U311 ( .A(n301), .B(n302), .C(n303), .Z(n332) );
  GTECH_OAI21 U312 ( .A(n333), .B(n334), .C(n335), .Z(n303) );
  GTECH_XNOR4 U313 ( .A(n299), .B(n305), .C(n297), .D(n298), .Z(n331) );
  GTECH_ADD_ABC U314 ( .A(n336), .B(n337), .C(n338), .COUT(n298) );
  GTECH_XNOR3 U315 ( .A(n339), .B(n340), .C(n341), .Z(n337) );
  GTECH_XOR2 U316 ( .A(n318), .B(n342), .Z(n297) );
  GTECH_AND2 U317 ( .A(I_b[6]), .B(I_a[0]), .Z(n342) );
  GTECH_XNOR3 U318 ( .A(n343), .B(n344), .C(n345), .Z(n318) );
  GTECH_NOT U319 ( .A(n314), .Z(n345) );
  GTECH_NAND3 U320 ( .A(I_b[4]), .B(I_a[1]), .C(n346), .Z(n314) );
  GTECH_NOT U321 ( .A(n313), .Z(n344) );
  GTECH_NAND2 U322 ( .A(I_b[5]), .B(I_a[1]), .Z(n313) );
  GTECH_NOT U323 ( .A(n312), .Z(n343) );
  GTECH_NAND2 U324 ( .A(I_b[4]), .B(I_a[2]), .Z(n312) );
  GTECH_NOT U325 ( .A(n300), .Z(n305) );
  GTECH_XNOR3 U326 ( .A(n322), .B(n324), .C(n319), .Z(n300) );
  GTECH_NOT U327 ( .A(n323), .Z(n319) );
  GTECH_OAI21 U328 ( .A(n347), .B(n348), .C(n349), .Z(n323) );
  GTECH_OAI21 U329 ( .A(n350), .B(n351), .C(n352), .Z(n349) );
  GTECH_NOT U330 ( .A(n353), .Z(n324) );
  GTECH_NAND2 U331 ( .A(I_b[3]), .B(I_a[3]), .Z(n353) );
  GTECH_NOT U332 ( .A(n320), .Z(n322) );
  GTECH_NAND2 U333 ( .A(I_b[2]), .B(I_a[4]), .Z(n320) );
  GTECH_NOT U334 ( .A(n354), .Z(n299) );
  GTECH_XNOR3 U335 ( .A(n306), .B(n307), .C(n327), .Z(n354) );
  GTECH_NOT U336 ( .A(n308), .Z(n327) );
  GTECH_OAI21 U337 ( .A(n355), .B(n356), .C(n357), .Z(n308) );
  GTECH_OAI21 U338 ( .A(n339), .B(n341), .C(n340), .Z(n357) );
  GTECH_NOT U339 ( .A(n358), .Z(n307) );
  GTECH_NAND2 U340 ( .A(I_a[5]), .B(I_b[1]), .Z(n358) );
  GTECH_NOT U341 ( .A(n328), .Z(n306) );
  GTECH_NAND2 U342 ( .A(I_a[6]), .B(I_b[0]), .Z(n328) );
  GTECH_XNOR3 U343 ( .A(n335), .B(n302), .C(n334), .Z(N145) );
  GTECH_NOT U344 ( .A(n301), .Z(n334) );
  GTECH_XOR2 U345 ( .A(n359), .B(n346), .Z(n301) );
  GTECH_NOT U346 ( .A(n360), .Z(n346) );
  GTECH_NAND2 U347 ( .A(I_b[5]), .B(I_a[0]), .Z(n360) );
  GTECH_NAND2 U348 ( .A(I_b[4]), .B(I_a[1]), .Z(n359) );
  GTECH_NOT U349 ( .A(n333), .Z(n302) );
  GTECH_XOR2 U350 ( .A(n361), .B(n336), .Z(n333) );
  GTECH_ADD_ABC U351 ( .A(n362), .B(n363), .C(n364), .COUT(n336) );
  GTECH_XNOR3 U352 ( .A(n365), .B(n366), .C(n367), .Z(n363) );
  GTECH_OA21 U353 ( .A(n368), .B(n369), .C(n370), .Z(n362) );
  GTECH_XNOR4 U354 ( .A(n340), .B(n355), .C(n338), .D(n339), .Z(n361) );
  GTECH_NOT U355 ( .A(n356), .Z(n339) );
  GTECH_NAND2 U356 ( .A(I_a[5]), .B(I_b[0]), .Z(n356) );
  GTECH_NOT U357 ( .A(n371), .Z(n338) );
  GTECH_XNOR3 U358 ( .A(n350), .B(n352), .C(n347), .Z(n371) );
  GTECH_NOT U359 ( .A(n351), .Z(n347) );
  GTECH_OAI21 U360 ( .A(n372), .B(n373), .C(n374), .Z(n351) );
  GTECH_NOT U361 ( .A(n375), .Z(n352) );
  GTECH_NAND2 U362 ( .A(I_b[3]), .B(I_a[2]), .Z(n375) );
  GTECH_NOT U363 ( .A(n348), .Z(n350) );
  GTECH_NAND2 U364 ( .A(I_b[2]), .B(I_a[3]), .Z(n348) );
  GTECH_NOT U365 ( .A(n341), .Z(n355) );
  GTECH_OAI21 U366 ( .A(n376), .B(n377), .C(n378), .Z(n341) );
  GTECH_OAI21 U367 ( .A(n365), .B(n367), .C(n366), .Z(n378) );
  GTECH_NOT U368 ( .A(n379), .Z(n340) );
  GTECH_NAND2 U369 ( .A(I_a[4]), .B(I_b[1]), .Z(n379) );
  GTECH_NOT U370 ( .A(n380), .Z(n335) );
  GTECH_NAND3 U371 ( .A(I_a[0]), .B(n381), .C(I_b[4]), .Z(n380) );
  GTECH_XOR2 U372 ( .A(n382), .B(n381), .Z(N144) );
  GTECH_XOR2 U373 ( .A(n383), .B(n384), .Z(n381) );
  GTECH_OA21 U374 ( .A(n368), .B(n369), .C(n370), .Z(n384) );
  GTECH_OAI21 U375 ( .A(n385), .B(n386), .C(n387), .Z(n370) );
  GTECH_XNOR4 U376 ( .A(n366), .B(n376), .C(n364), .D(n365), .Z(n383) );
  GTECH_NOT U377 ( .A(n377), .Z(n365) );
  GTECH_NAND2 U378 ( .A(I_a[4]), .B(I_b[0]), .Z(n377) );
  GTECH_XNOR3 U379 ( .A(n388), .B(n389), .C(n390), .Z(n364) );
  GTECH_NOT U380 ( .A(n374), .Z(n390) );
  GTECH_NAND3 U381 ( .A(I_b[2]), .B(I_a[1]), .C(n391), .Z(n374) );
  GTECH_NOT U382 ( .A(n373), .Z(n389) );
  GTECH_NAND2 U383 ( .A(I_b[3]), .B(I_a[1]), .Z(n373) );
  GTECH_NOT U384 ( .A(n372), .Z(n388) );
  GTECH_NAND2 U385 ( .A(I_b[2]), .B(I_a[2]), .Z(n372) );
  GTECH_NOT U386 ( .A(n367), .Z(n376) );
  GTECH_OAI21 U387 ( .A(n392), .B(n393), .C(n394), .Z(n367) );
  GTECH_OAI21 U388 ( .A(n395), .B(n396), .C(n397), .Z(n394) );
  GTECH_NOT U389 ( .A(n398), .Z(n366) );
  GTECH_NAND2 U390 ( .A(I_a[3]), .B(I_b[1]), .Z(n398) );
  GTECH_AND2 U391 ( .A(I_b[4]), .B(I_a[0]), .Z(n382) );
  GTECH_XNOR3 U392 ( .A(n387), .B(n369), .C(n386), .Z(N143) );
  GTECH_NOT U393 ( .A(n368), .Z(n386) );
  GTECH_XOR2 U394 ( .A(n399), .B(n391), .Z(n368) );
  GTECH_NOT U395 ( .A(n400), .Z(n391) );
  GTECH_NAND2 U396 ( .A(I_b[3]), .B(I_a[0]), .Z(n400) );
  GTECH_NAND2 U397 ( .A(I_b[2]), .B(I_a[1]), .Z(n399) );
  GTECH_NOT U398 ( .A(n385), .Z(n369) );
  GTECH_XNOR3 U399 ( .A(n395), .B(n397), .C(n392), .Z(n385) );
  GTECH_NOT U400 ( .A(n396), .Z(n392) );
  GTECH_OAI21 U401 ( .A(n401), .B(n402), .C(n403), .Z(n396) );
  GTECH_NOT U402 ( .A(n404), .Z(n397) );
  GTECH_NAND2 U403 ( .A(I_b[1]), .B(I_a[2]), .Z(n404) );
  GTECH_NOT U404 ( .A(n393), .Z(n395) );
  GTECH_NAND2 U405 ( .A(I_b[0]), .B(I_a[3]), .Z(n393) );
  GTECH_NOT U406 ( .A(n405), .Z(n387) );
  GTECH_NAND3 U407 ( .A(I_a[0]), .B(n406), .C(I_b[2]), .Z(n405) );
  GTECH_XOR2 U408 ( .A(n407), .B(n406), .Z(N142) );
  GTECH_NOT U409 ( .A(n408), .Z(n406) );
  GTECH_XNOR3 U410 ( .A(n409), .B(n410), .C(n411), .Z(n408) );
  GTECH_NOT U411 ( .A(n403), .Z(n411) );
  GTECH_NAND3 U412 ( .A(n412), .B(I_b[0]), .C(I_a[1]), .Z(n403) );
  GTECH_NOT U413 ( .A(n401), .Z(n410) );
  GTECH_NAND2 U414 ( .A(I_a[1]), .B(I_b[1]), .Z(n401) );
  GTECH_NOT U415 ( .A(n402), .Z(n409) );
  GTECH_NAND2 U416 ( .A(I_b[0]), .B(I_a[2]), .Z(n402) );
  GTECH_AND2 U417 ( .A(I_b[2]), .B(I_a[0]), .Z(n407) );
  GTECH_XOR2 U418 ( .A(n412), .B(n413), .Z(N141) );
  GTECH_AND2 U419 ( .A(I_a[1]), .B(I_b[0]), .Z(n413) );
  GTECH_NOT U420 ( .A(n414), .Z(n412) );
  GTECH_NAND2 U421 ( .A(I_a[0]), .B(I_b[1]), .Z(n414) );
  GTECH_AND2 U422 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

