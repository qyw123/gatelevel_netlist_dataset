
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374;

  GTECH_MUX2 U131 ( .A(n270), .B(n271), .S(n272), .Z(sum[9]) );
  GTECH_OA21 U132 ( .A(n273), .B(n274), .C(n275), .Z(n272) );
  GTECH_NOT U133 ( .A(n276), .Z(n274) );
  GTECH_XOR2 U134 ( .A(b[9]), .B(a[9]), .Z(n271) );
  GTECH_OR_NOT U135 ( .A(n277), .B(n278), .Z(n270) );
  GTECH_XNOR2 U136 ( .A(n279), .B(n276), .Z(sum[8]) );
  GTECH_MUX2 U137 ( .A(n280), .B(n281), .S(n282), .Z(sum[7]) );
  GTECH_XNOR2 U138 ( .A(n283), .B(n284), .Z(n281) );
  GTECH_XOR2 U139 ( .A(n283), .B(n285), .Z(n280) );
  GTECH_AND_NOT U140 ( .A(n286), .B(n287), .Z(n285) );
  GTECH_OAI21 U141 ( .A(b[6]), .B(a[6]), .C(n288), .Z(n286) );
  GTECH_XNOR2 U142 ( .A(a[7]), .B(b[7]), .Z(n283) );
  GTECH_AO21 U143 ( .A(n289), .B(n287), .C(n290), .Z(sum[6]) );
  GTECH_NOT U144 ( .A(n291), .Z(n290) );
  GTECH_MUX2 U145 ( .A(n292), .B(n293), .S(b[6]), .Z(n291) );
  GTECH_OR2 U146 ( .A(n289), .B(a[6]), .Z(n293) );
  GTECH_XNOR2 U147 ( .A(a[6]), .B(n289), .Z(n292) );
  GTECH_AO21 U148 ( .A(n294), .B(n282), .C(n288), .Z(n289) );
  GTECH_OA21 U149 ( .A(n295), .B(n296), .C(n297), .Z(n288) );
  GTECH_MUX2 U150 ( .A(n298), .B(n299), .S(n300), .Z(sum[5]) );
  GTECH_AND_NOT U151 ( .A(n297), .B(n296), .Z(n300) );
  GTECH_OAI21 U152 ( .A(n295), .B(n282), .C(n301), .Z(n299) );
  GTECH_AO21 U153 ( .A(n301), .B(n282), .C(n295), .Z(n298) );
  GTECH_XOR2 U154 ( .A(n282), .B(n302), .Z(sum[4]) );
  GTECH_MUX2 U155 ( .A(n303), .B(n304), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U156 ( .A(n305), .B(n306), .Z(n304) );
  GTECH_XNOR2 U157 ( .A(n305), .B(n307), .Z(n303) );
  GTECH_AND_NOT U158 ( .A(n308), .B(n309), .Z(n307) );
  GTECH_AO21 U159 ( .A(n310), .B(n311), .C(n312), .Z(n308) );
  GTECH_XOR2 U160 ( .A(a[3]), .B(b[3]), .Z(n305) );
  GTECH_MUX2 U161 ( .A(n313), .B(n314), .S(cin), .Z(sum[2]) );
  GTECH_MUX2 U162 ( .A(n315), .B(n316), .S(n317), .Z(n314) );
  GTECH_MUX2 U163 ( .A(n315), .B(n316), .S(n312), .Z(n313) );
  GTECH_OAI21 U164 ( .A(n318), .B(n319), .C(n320), .Z(n312) );
  GTECH_XOR2 U165 ( .A(a[2]), .B(b[2]), .Z(n316) );
  GTECH_AO21 U166 ( .A(n310), .B(n311), .C(n309), .Z(n315) );
  GTECH_MUX2 U167 ( .A(n321), .B(n322), .S(n323), .Z(sum[1]) );
  GTECH_AND_NOT U168 ( .A(n320), .B(n319), .Z(n323) );
  GTECH_OAI21 U169 ( .A(cin), .B(n318), .C(n324), .Z(n322) );
  GTECH_AO21 U170 ( .A(n324), .B(cin), .C(n318), .Z(n321) );
  GTECH_MUX2 U171 ( .A(n325), .B(n326), .S(n327), .Z(sum[15]) );
  GTECH_XOR2 U172 ( .A(n328), .B(n329), .Z(n326) );
  GTECH_OA21 U173 ( .A(n330), .B(n331), .C(n332), .Z(n329) );
  GTECH_XNOR2 U174 ( .A(n328), .B(n333), .Z(n325) );
  GTECH_XNOR2 U175 ( .A(a[15]), .B(b[15]), .Z(n328) );
  GTECH_MUX2 U176 ( .A(n334), .B(n335), .S(n336), .Z(sum[14]) );
  GTECH_OA21 U177 ( .A(n327), .B(n337), .C(n331), .Z(n336) );
  GTECH_OAI22 U178 ( .A(b[13]), .B(a[13]), .C(n338), .D(n339), .Z(n331) );
  GTECH_XOR2 U179 ( .A(b[14]), .B(a[14]), .Z(n335) );
  GTECH_OR_NOT U180 ( .A(n330), .B(n332), .Z(n334) );
  GTECH_MUX2 U181 ( .A(n340), .B(n341), .S(n327), .Z(sum[13]) );
  GTECH_MUX2 U182 ( .A(n342), .B(n343), .S(n339), .Z(n341) );
  GTECH_MUX2 U183 ( .A(n342), .B(n343), .S(n344), .Z(n340) );
  GTECH_OAI21 U184 ( .A(a[13]), .B(b[13]), .C(n345), .Z(n343) );
  GTECH_NOT U185 ( .A(n338), .Z(n345) );
  GTECH_XNOR2 U186 ( .A(n346), .B(b[13]), .Z(n342) );
  GTECH_NOT U187 ( .A(a[13]), .Z(n346) );
  GTECH_XNOR2 U188 ( .A(n347), .B(n327), .Z(sum[12]) );
  GTECH_MUX2 U189 ( .A(n348), .B(n349), .S(n276), .Z(sum[11]) );
  GTECH_XNOR2 U190 ( .A(n350), .B(n351), .Z(n349) );
  GTECH_XOR2 U191 ( .A(n350), .B(n352), .Z(n348) );
  GTECH_AND_NOT U192 ( .A(n353), .B(n354), .Z(n352) );
  GTECH_OAI21 U193 ( .A(b[10]), .B(a[10]), .C(n355), .Z(n353) );
  GTECH_XNOR2 U194 ( .A(a[11]), .B(b[11]), .Z(n350) );
  GTECH_AO21 U195 ( .A(n356), .B(n354), .C(n357), .Z(sum[10]) );
  GTECH_NOT U196 ( .A(n358), .Z(n357) );
  GTECH_MUX2 U197 ( .A(n359), .B(n360), .S(b[10]), .Z(n358) );
  GTECH_OR2 U198 ( .A(n356), .B(a[10]), .Z(n360) );
  GTECH_XNOR2 U199 ( .A(a[10]), .B(n356), .Z(n359) );
  GTECH_AO21 U200 ( .A(n361), .B(n276), .C(n355), .Z(n356) );
  GTECH_OAI21 U201 ( .A(n277), .B(n275), .C(n278), .Z(n355) );
  GTECH_XOR2 U202 ( .A(cin), .B(n362), .Z(sum[0]) );
  GTECH_MUX2 U203 ( .A(n363), .B(n347), .S(n327), .Z(cout) );
  GTECH_MUX2 U204 ( .A(n279), .B(n364), .S(n276), .Z(n327) );
  GTECH_MUX2 U205 ( .A(n302), .B(n365), .S(n282), .Z(n276) );
  GTECH_MUX2 U206 ( .A(n362), .B(n366), .S(cin), .Z(n282) );
  GTECH_OA21 U207 ( .A(a[3]), .B(n306), .C(n367), .Z(n366) );
  GTECH_AO21 U208 ( .A(n306), .B(a[3]), .C(b[3]), .Z(n367) );
  GTECH_OR_NOT U209 ( .A(n309), .B(n368), .Z(n306) );
  GTECH_AO21 U210 ( .A(n311), .B(n310), .C(n317), .Z(n368) );
  GTECH_OAI21 U211 ( .A(n319), .B(n324), .C(n320), .Z(n317) );
  GTECH_OR2 U212 ( .A(b[1]), .B(a[1]), .Z(n320) );
  GTECH_AND2 U213 ( .A(b[1]), .B(a[1]), .Z(n319) );
  GTECH_NOT U214 ( .A(b[2]), .Z(n310) );
  GTECH_NOT U215 ( .A(a[2]), .Z(n311) );
  GTECH_AND2 U216 ( .A(b[2]), .B(a[2]), .Z(n309) );
  GTECH_AND_NOT U217 ( .A(n324), .B(n318), .Z(n362) );
  GTECH_AND2 U218 ( .A(a[0]), .B(b[0]), .Z(n318) );
  GTECH_OR2 U219 ( .A(b[0]), .B(a[0]), .Z(n324) );
  GTECH_AO21 U220 ( .A(n284), .B(a[7]), .C(n369), .Z(n365) );
  GTECH_OA21 U221 ( .A(a[7]), .B(n284), .C(b[7]), .Z(n369) );
  GTECH_OR_NOT U222 ( .A(n287), .B(n370), .Z(n284) );
  GTECH_OAI21 U223 ( .A(a[6]), .B(b[6]), .C(n294), .Z(n370) );
  GTECH_OA21 U224 ( .A(n296), .B(n301), .C(n297), .Z(n294) );
  GTECH_OR2 U225 ( .A(b[5]), .B(a[5]), .Z(n297) );
  GTECH_AND2 U226 ( .A(a[5]), .B(b[5]), .Z(n296) );
  GTECH_AND2 U227 ( .A(b[6]), .B(a[6]), .Z(n287) );
  GTECH_AND_NOT U228 ( .A(n301), .B(n295), .Z(n302) );
  GTECH_AND2 U229 ( .A(b[4]), .B(a[4]), .Z(n295) );
  GTECH_OR2 U230 ( .A(a[4]), .B(b[4]), .Z(n301) );
  GTECH_NOT U231 ( .A(n371), .Z(n364) );
  GTECH_AO21 U232 ( .A(n351), .B(a[11]), .C(n372), .Z(n371) );
  GTECH_OA21 U233 ( .A(a[11]), .B(n351), .C(b[11]), .Z(n372) );
  GTECH_OR_NOT U234 ( .A(n354), .B(n373), .Z(n351) );
  GTECH_OAI21 U235 ( .A(a[10]), .B(b[10]), .C(n361), .Z(n373) );
  GTECH_OAI21 U236 ( .A(n277), .B(n273), .C(n278), .Z(n361) );
  GTECH_NAND2 U237 ( .A(b[9]), .B(a[9]), .Z(n278) );
  GTECH_NOR2 U238 ( .A(b[9]), .B(a[9]), .Z(n277) );
  GTECH_AND2 U239 ( .A(b[10]), .B(a[10]), .Z(n354) );
  GTECH_OR_NOT U240 ( .A(n273), .B(n275), .Z(n279) );
  GTECH_NAND2 U241 ( .A(a[8]), .B(b[8]), .Z(n275) );
  GTECH_NOR2 U242 ( .A(b[8]), .B(a[8]), .Z(n273) );
  GTECH_AND_NOT U243 ( .A(n344), .B(n339), .Z(n347) );
  GTECH_AND2 U244 ( .A(b[12]), .B(a[12]), .Z(n339) );
  GTECH_AO21 U245 ( .A(n333), .B(a[15]), .C(n374), .Z(n363) );
  GTECH_OA21 U246 ( .A(a[15]), .B(n333), .C(b[15]), .Z(n374) );
  GTECH_OAI21 U247 ( .A(n330), .B(n337), .C(n332), .Z(n333) );
  GTECH_NAND2 U248 ( .A(a[14]), .B(b[14]), .Z(n332) );
  GTECH_OAI22 U249 ( .A(b[13]), .B(a[13]), .C(n338), .D(n344), .Z(n337) );
  GTECH_OR2 U250 ( .A(b[12]), .B(a[12]), .Z(n344) );
  GTECH_AND2 U251 ( .A(b[13]), .B(a[13]), .Z(n338) );
  GTECH_NOR2 U252 ( .A(a[14]), .B(b[14]), .Z(n330) );
endmodule

