
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_OR_NOT U83 ( .A(n97), .B(n93), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n98), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n98) );
  GTECH_OAI21 U86 ( .A(n99), .B(n100), .C(n101), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  GTECH_NOT U88 ( .A(n103), .Z(n99) );
  GTECH_OR_NOT U89 ( .A(n105), .B(I_b[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n106), .Z(n84) );
  GTECH_OR_NOT U91 ( .A(n107), .B(n108), .Z(n106) );
  GTECH_XOR2 U92 ( .A(n109), .B(n108), .Z(N153) );
  GTECH_NOT U93 ( .A(n110), .Z(n108) );
  GTECH_XOR3 U94 ( .A(n97), .B(n93), .C(n95), .Z(n110) );
  GTECH_XOR3 U95 ( .A(n102), .B(n104), .C(n103), .Z(n95) );
  GTECH_OAI21 U96 ( .A(n111), .B(n112), .C(n113), .Z(n103) );
  GTECH_OAI21 U97 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_NOT U98 ( .A(n115), .Z(n111) );
  GTECH_NOT U99 ( .A(n117), .Z(n104) );
  GTECH_OR_NOT U100 ( .A(n118), .B(I_b[7]), .Z(n117) );
  GTECH_NOT U101 ( .A(n100), .Z(n102) );
  GTECH_OR_NOT U102 ( .A(n119), .B(I_a[7]), .Z(n100) );
  GTECH_NOT U103 ( .A(I_b[6]), .Z(n119) );
  GTECH_ADD_ABC U104 ( .A(n120), .B(n121), .C(n122), .COUT(n93) );
  GTECH_NOT U105 ( .A(n123), .Z(n122) );
  GTECH_XOR2 U106 ( .A(n124), .B(n125), .Z(n121) );
  GTECH_AND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n125) );
  GTECH_NOT U108 ( .A(n94), .Z(n97) );
  GTECH_OR_NOT U109 ( .A(n124), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U110 ( .A(n107), .Z(n109) );
  GTECH_OR_NOT U111 ( .A(n126), .B(n127), .Z(n107) );
  GTECH_XOR2 U112 ( .A(n126), .B(n128), .Z(N152) );
  GTECH_NOT U113 ( .A(n127), .Z(n128) );
  GTECH_XOR4 U114 ( .A(n129), .B(n124), .C(n120), .D(n123), .Z(n127) );
  GTECH_XOR3 U115 ( .A(n114), .B(n116), .C(n115), .Z(n123) );
  GTECH_OAI21 U116 ( .A(n130), .B(n131), .C(n132), .Z(n115) );
  GTECH_OAI21 U117 ( .A(n133), .B(n134), .C(n135), .Z(n132) );
  GTECH_NOT U118 ( .A(n134), .Z(n130) );
  GTECH_NOT U119 ( .A(n136), .Z(n116) );
  GTECH_OR_NOT U120 ( .A(n137), .B(I_b[7]), .Z(n136) );
  GTECH_NOT U121 ( .A(n112), .Z(n114) );
  GTECH_OR_NOT U122 ( .A(n118), .B(I_b[6]), .Z(n112) );
  GTECH_NOT U123 ( .A(I_a[6]), .Z(n118) );
  GTECH_ADD_ABC U124 ( .A(n138), .B(n139), .C(n140), .COUT(n120) );
  GTECH_NOT U125 ( .A(n141), .Z(n140) );
  GTECH_XOR3 U126 ( .A(n142), .B(n143), .C(n144), .Z(n139) );
  GTECH_NOT U127 ( .A(n145), .Z(n142) );
  GTECH_OA22 U128 ( .A(n144), .B(n145), .C(n146), .D(n147), .Z(n124) );
  GTECH_AND_NOT U129 ( .A(n145), .B(n148), .Z(n146) );
  GTECH_NOT U130 ( .A(n148), .Z(n144) );
  GTECH_AND2 U131 ( .A(I_b[5]), .B(I_a[7]), .Z(n129) );
  GTECH_ADD_ABC U132 ( .A(n149), .B(n150), .C(n151), .COUT(n126) );
  GTECH_NOT U133 ( .A(n152), .Z(n151) );
  GTECH_OA22 U134 ( .A(n153), .B(n105), .C(n154), .D(n155), .Z(n150) );
  GTECH_OA22 U135 ( .A(n156), .B(n157), .C(n158), .D(n159), .Z(n149) );
  GTECH_AND2 U136 ( .A(n158), .B(n159), .Z(n156) );
  GTECH_XOR3 U137 ( .A(n160), .B(n152), .C(n161), .Z(N151) );
  GTECH_AOI2N2 U138 ( .A(n162), .B(n163), .C(n158), .D(n159), .Z(n161) );
  GTECH_OR_NOT U139 ( .A(n164), .B(n159), .Z(n163) );
  GTECH_XOR2 U140 ( .A(n165), .B(n138), .Z(n152) );
  GTECH_ADD_ABC U141 ( .A(n166), .B(n167), .C(n168), .COUT(n138) );
  GTECH_NOT U142 ( .A(n169), .Z(n168) );
  GTECH_XOR3 U143 ( .A(n170), .B(n171), .C(n172), .Z(n167) );
  GTECH_XOR4 U144 ( .A(n143), .B(n148), .C(n145), .D(n141), .Z(n165) );
  GTECH_XOR3 U145 ( .A(n133), .B(n135), .C(n134), .Z(n141) );
  GTECH_OAI21 U146 ( .A(n173), .B(n174), .C(n175), .Z(n134) );
  GTECH_OAI21 U147 ( .A(n176), .B(n177), .C(n178), .Z(n175) );
  GTECH_NOT U148 ( .A(n177), .Z(n173) );
  GTECH_NOT U149 ( .A(n179), .Z(n135) );
  GTECH_OR_NOT U150 ( .A(n180), .B(I_b[7]), .Z(n179) );
  GTECH_NOT U151 ( .A(n131), .Z(n133) );
  GTECH_OR_NOT U152 ( .A(n137), .B(I_b[6]), .Z(n131) );
  GTECH_NOT U153 ( .A(I_a[5]), .Z(n137) );
  GTECH_OR_NOT U154 ( .A(n181), .B(I_a[7]), .Z(n145) );
  GTECH_OAI21 U155 ( .A(n172), .B(n182), .C(n183), .Z(n148) );
  GTECH_OAI21 U156 ( .A(n170), .B(n184), .C(n171), .Z(n183) );
  GTECH_NOT U157 ( .A(n182), .Z(n170) );
  GTECH_NOT U158 ( .A(n184), .Z(n172) );
  GTECH_NOT U159 ( .A(n147), .Z(n143) );
  GTECH_OR_NOT U160 ( .A(n185), .B(I_a[6]), .Z(n147) );
  GTECH_OA22 U161 ( .A(n153), .B(n105), .C(n154), .D(n155), .Z(n160) );
  GTECH_NOT U162 ( .A(n186), .Z(n155) );
  GTECH_NOT U163 ( .A(I_a[7]), .Z(n105) );
  GTECH_XOR3 U164 ( .A(n158), .B(n187), .C(n157), .Z(N150) );
  GTECH_NOT U165 ( .A(n162), .Z(n157) );
  GTECH_XOR2 U166 ( .A(n188), .B(n166), .Z(n162) );
  GTECH_ADD_ABC U167 ( .A(n189), .B(n190), .C(n191), .COUT(n166) );
  GTECH_NOT U168 ( .A(n192), .Z(n191) );
  GTECH_XOR3 U169 ( .A(n193), .B(n194), .C(n195), .Z(n190) );
  GTECH_XOR4 U170 ( .A(n171), .B(n184), .C(n182), .D(n169), .Z(n188) );
  GTECH_XOR3 U171 ( .A(n176), .B(n178), .C(n177), .Z(n169) );
  GTECH_OAI21 U172 ( .A(n196), .B(n197), .C(n198), .Z(n177) );
  GTECH_OAI21 U173 ( .A(n199), .B(n200), .C(n201), .Z(n198) );
  GTECH_NOT U174 ( .A(n200), .Z(n196) );
  GTECH_NOT U175 ( .A(n202), .Z(n178) );
  GTECH_OR_NOT U176 ( .A(n203), .B(I_b[7]), .Z(n202) );
  GTECH_NOT U177 ( .A(n174), .Z(n176) );
  GTECH_OR_NOT U178 ( .A(n180), .B(I_b[6]), .Z(n174) );
  GTECH_OR_NOT U179 ( .A(n181), .B(I_a[6]), .Z(n182) );
  GTECH_OAI21 U180 ( .A(n195), .B(n204), .C(n205), .Z(n184) );
  GTECH_OAI21 U181 ( .A(n193), .B(n206), .C(n194), .Z(n205) );
  GTECH_NOT U182 ( .A(n204), .Z(n193) );
  GTECH_NOT U183 ( .A(n206), .Z(n195) );
  GTECH_NOT U184 ( .A(n207), .Z(n171) );
  GTECH_OR_NOT U185 ( .A(n185), .B(I_a[5]), .Z(n207) );
  GTECH_NOT U186 ( .A(I_b[5]), .Z(n185) );
  GTECH_NOT U187 ( .A(n159), .Z(n187) );
  GTECH_XOR2 U188 ( .A(n186), .B(n154), .Z(n159) );
  GTECH_AOI2N2 U189 ( .A(n208), .B(n209), .C(n210), .D(n211), .Z(n154) );
  GTECH_OR_NOT U190 ( .A(n212), .B(n210), .Z(n209) );
  GTECH_XOR2 U191 ( .A(n213), .B(n153), .Z(n186) );
  GTECH_AND2 U192 ( .A(n214), .B(n215), .Z(n153) );
  GTECH_OR_NOT U193 ( .A(n216), .B(n217), .Z(n215) );
  GTECH_OAI21 U194 ( .A(n218), .B(n217), .C(n219), .Z(n214) );
  GTECH_OR_NOT U195 ( .A(n220), .B(I_a[7]), .Z(n213) );
  GTECH_NOT U196 ( .A(n164), .Z(n158) );
  GTECH_OAI2N2 U197 ( .A(n221), .B(n222), .C(n223), .D(n224), .Z(n164) );
  GTECH_OR_NOT U198 ( .A(n225), .B(n221), .Z(n224) );
  GTECH_XOR3 U199 ( .A(n221), .B(n225), .C(n226), .Z(N149) );
  GTECH_NOT U200 ( .A(n223), .Z(n226) );
  GTECH_XOR2 U201 ( .A(n227), .B(n189), .Z(n223) );
  GTECH_ADD_ABC U202 ( .A(n228), .B(n229), .C(n230), .COUT(n189) );
  GTECH_XOR3 U203 ( .A(n231), .B(n232), .C(n233), .Z(n229) );
  GTECH_OA22 U204 ( .A(n234), .B(n235), .C(n236), .D(n237), .Z(n228) );
  GTECH_AND2 U205 ( .A(n236), .B(n237), .Z(n234) );
  GTECH_XOR4 U206 ( .A(n194), .B(n206), .C(n204), .D(n192), .Z(n227) );
  GTECH_XOR3 U207 ( .A(n199), .B(n201), .C(n200), .Z(n192) );
  GTECH_OAI21 U208 ( .A(n238), .B(n239), .C(n240), .Z(n200) );
  GTECH_NOT U209 ( .A(n241), .Z(n201) );
  GTECH_OR_NOT U210 ( .A(n242), .B(I_b[7]), .Z(n241) );
  GTECH_NOT U211 ( .A(n197), .Z(n199) );
  GTECH_OR_NOT U212 ( .A(n203), .B(I_b[6]), .Z(n197) );
  GTECH_OR_NOT U213 ( .A(n181), .B(I_a[5]), .Z(n204) );
  GTECH_NOT U214 ( .A(I_b[4]), .Z(n181) );
  GTECH_OAI21 U215 ( .A(n233), .B(n243), .C(n244), .Z(n206) );
  GTECH_OAI21 U216 ( .A(n231), .B(n245), .C(n232), .Z(n244) );
  GTECH_NOT U217 ( .A(n243), .Z(n231) );
  GTECH_NOT U218 ( .A(n245), .Z(n233) );
  GTECH_NOT U219 ( .A(n246), .Z(n194) );
  GTECH_OR_NOT U220 ( .A(n180), .B(I_b[5]), .Z(n246) );
  GTECH_NOT U221 ( .A(n222), .Z(n225) );
  GTECH_XOR3 U222 ( .A(n212), .B(n210), .C(n208), .Z(n222) );
  GTECH_XOR3 U223 ( .A(n218), .B(n219), .C(n217), .Z(n208) );
  GTECH_OAI21 U224 ( .A(n247), .B(n248), .C(n249), .Z(n217) );
  GTECH_OAI21 U225 ( .A(n250), .B(n251), .C(n252), .Z(n249) );
  GTECH_NOT U226 ( .A(n251), .Z(n247) );
  GTECH_NOT U227 ( .A(n253), .Z(n219) );
  GTECH_OR_NOT U228 ( .A(n220), .B(I_a[6]), .Z(n253) );
  GTECH_NOT U229 ( .A(n216), .Z(n218) );
  GTECH_OR_NOT U230 ( .A(n254), .B(I_a[7]), .Z(n216) );
  GTECH_ADD_ABC U231 ( .A(n255), .B(n256), .C(n257), .COUT(n210) );
  GTECH_XOR2 U232 ( .A(n258), .B(n259), .Z(n256) );
  GTECH_AND2 U233 ( .A(I_a[7]), .B(I_b[1]), .Z(n259) );
  GTECH_NOT U234 ( .A(n211), .Z(n212) );
  GTECH_OR_NOT U235 ( .A(n258), .B(I_a[7]), .Z(n211) );
  GTECH_ADD_ABC U236 ( .A(n260), .B(n261), .C(n262), .COUT(n221) );
  GTECH_XOR3 U237 ( .A(n255), .B(n263), .C(n257), .Z(n261) );
  GTECH_NOT U238 ( .A(n264), .Z(n257) );
  GTECH_XOR2 U239 ( .A(n260), .B(n265), .Z(N148) );
  GTECH_XOR4 U240 ( .A(n263), .B(n264), .C(n262), .D(n255), .Z(n265) );
  GTECH_ADD_ABC U241 ( .A(n266), .B(n267), .C(n268), .COUT(n255) );
  GTECH_XOR3 U242 ( .A(n269), .B(n270), .C(n271), .Z(n267) );
  GTECH_XOR2 U243 ( .A(n272), .B(n273), .Z(n262) );
  GTECH_OA22 U244 ( .A(n236), .B(n237), .C(n274), .D(n235), .Z(n273) );
  GTECH_AND_NOT U245 ( .A(n236), .B(n275), .Z(n274) );
  GTECH_XOR4 U246 ( .A(n232), .B(n245), .C(n243), .D(n230), .Z(n272) );
  GTECH_XOR3 U247 ( .A(n276), .B(n277), .C(n240), .Z(n230) );
  GTECH_NAND3 U248 ( .A(I_b[6]), .B(I_a[1]), .C(n278), .Z(n240) );
  GTECH_NOT U249 ( .A(n239), .Z(n277) );
  GTECH_OR_NOT U250 ( .A(n279), .B(I_b[7]), .Z(n239) );
  GTECH_NOT U251 ( .A(n238), .Z(n276) );
  GTECH_OR_NOT U252 ( .A(n242), .B(I_b[6]), .Z(n238) );
  GTECH_OR_NOT U253 ( .A(n180), .B(I_b[4]), .Z(n243) );
  GTECH_OAI21 U254 ( .A(n280), .B(n281), .C(n282), .Z(n245) );
  GTECH_OAI21 U255 ( .A(n283), .B(n284), .C(n285), .Z(n282) );
  GTECH_NOT U256 ( .A(n284), .Z(n280) );
  GTECH_NOT U257 ( .A(n286), .Z(n232) );
  GTECH_OR_NOT U258 ( .A(n203), .B(I_b[5]), .Z(n286) );
  GTECH_XOR3 U259 ( .A(n250), .B(n252), .C(n251), .Z(n264) );
  GTECH_OAI21 U260 ( .A(n287), .B(n288), .C(n289), .Z(n251) );
  GTECH_OAI21 U261 ( .A(n290), .B(n291), .C(n292), .Z(n289) );
  GTECH_NOT U262 ( .A(n291), .Z(n287) );
  GTECH_NOT U263 ( .A(n293), .Z(n252) );
  GTECH_OR_NOT U264 ( .A(n220), .B(I_a[5]), .Z(n293) );
  GTECH_NOT U265 ( .A(I_b[3]), .Z(n220) );
  GTECH_NOT U266 ( .A(n248), .Z(n250) );
  GTECH_OR_NOT U267 ( .A(n254), .B(I_a[6]), .Z(n248) );
  GTECH_XOR2 U268 ( .A(n294), .B(n258), .Z(n263) );
  GTECH_OA22 U269 ( .A(n271), .B(n295), .C(n296), .D(n297), .Z(n258) );
  GTECH_AND_NOT U270 ( .A(n295), .B(n298), .Z(n296) );
  GTECH_NOT U271 ( .A(n298), .Z(n271) );
  GTECH_AND2 U272 ( .A(I_b[1]), .B(I_a[7]), .Z(n294) );
  GTECH_ADD_ABC U273 ( .A(n299), .B(n300), .C(n301), .COUT(n260) );
  GTECH_NOT U274 ( .A(n302), .Z(n301) );
  GTECH_XOR3 U275 ( .A(n266), .B(n303), .C(n268), .Z(n300) );
  GTECH_NOT U276 ( .A(n304), .Z(n268) );
  GTECH_NOT U277 ( .A(n305), .Z(n303) );
  GTECH_XOR2 U278 ( .A(n306), .B(n299), .Z(N147) );
  GTECH_ADD_ABC U279 ( .A(n307), .B(n308), .C(n309), .COUT(n299) );
  GTECH_XOR3 U280 ( .A(n310), .B(n311), .C(n312), .Z(n308) );
  GTECH_OA22 U281 ( .A(n313), .B(n314), .C(n315), .D(n316), .Z(n307) );
  GTECH_AND2 U282 ( .A(n315), .B(n316), .Z(n313) );
  GTECH_XOR4 U283 ( .A(n304), .B(n266), .C(n305), .D(n302), .Z(n306) );
  GTECH_XOR3 U284 ( .A(n317), .B(n237), .C(n236), .Z(n302) );
  GTECH_XOR2 U285 ( .A(n318), .B(n278), .Z(n236) );
  GTECH_NOT U286 ( .A(n319), .Z(n278) );
  GTECH_OR_NOT U287 ( .A(n320), .B(I_b[7]), .Z(n319) );
  GTECH_OR_NOT U288 ( .A(n279), .B(I_b[6]), .Z(n318) );
  GTECH_NOT U289 ( .A(n275), .Z(n237) );
  GTECH_XOR3 U290 ( .A(n283), .B(n285), .C(n284), .Z(n275) );
  GTECH_OAI21 U291 ( .A(n321), .B(n322), .C(n323), .Z(n284) );
  GTECH_NOT U292 ( .A(n324), .Z(n285) );
  GTECH_OR_NOT U293 ( .A(n242), .B(I_b[5]), .Z(n324) );
  GTECH_NOT U294 ( .A(n281), .Z(n283) );
  GTECH_OR_NOT U295 ( .A(n203), .B(I_b[4]), .Z(n281) );
  GTECH_NOT U296 ( .A(n235), .Z(n317) );
  GTECH_NAND3 U297 ( .A(I_a[0]), .B(n325), .C(I_b[6]), .Z(n235) );
  GTECH_NOT U298 ( .A(n326), .Z(n325) );
  GTECH_XOR3 U299 ( .A(n269), .B(n270), .C(n298), .Z(n305) );
  GTECH_OAI21 U300 ( .A(n327), .B(n328), .C(n329), .Z(n298) );
  GTECH_OAI21 U301 ( .A(n330), .B(n331), .C(n332), .Z(n329) );
  GTECH_NOT U302 ( .A(n297), .Z(n270) );
  GTECH_OR_NOT U303 ( .A(n333), .B(I_a[6]), .Z(n297) );
  GTECH_NOT U304 ( .A(n295), .Z(n269) );
  GTECH_OR_NOT U305 ( .A(n334), .B(I_a[7]), .Z(n295) );
  GTECH_ADD_ABC U306 ( .A(n310), .B(n335), .C(n312), .COUT(n266) );
  GTECH_NOT U307 ( .A(n336), .Z(n312) );
  GTECH_XOR3 U308 ( .A(n330), .B(n332), .C(n327), .Z(n335) );
  GTECH_NOT U309 ( .A(n331), .Z(n327) );
  GTECH_XOR3 U310 ( .A(n290), .B(n292), .C(n291), .Z(n304) );
  GTECH_OAI21 U311 ( .A(n337), .B(n338), .C(n339), .Z(n291) );
  GTECH_OAI21 U312 ( .A(n340), .B(n341), .C(n342), .Z(n339) );
  GTECH_NOT U313 ( .A(n341), .Z(n337) );
  GTECH_NOT U314 ( .A(n343), .Z(n292) );
  GTECH_OR_NOT U315 ( .A(n180), .B(I_b[3]), .Z(n343) );
  GTECH_NOT U316 ( .A(n288), .Z(n290) );
  GTECH_OR_NOT U317 ( .A(n254), .B(I_a[5]), .Z(n288) );
  GTECH_NOT U318 ( .A(I_b[2]), .Z(n254) );
  GTECH_XOR2 U319 ( .A(n344), .B(n345), .Z(N146) );
  GTECH_XOR4 U320 ( .A(n311), .B(n336), .C(n309), .D(n310), .Z(n345) );
  GTECH_ADD_ABC U321 ( .A(n346), .B(n347), .C(n348), .COUT(n310) );
  GTECH_NOT U322 ( .A(n349), .Z(n348) );
  GTECH_XOR3 U323 ( .A(n350), .B(n351), .C(n352), .Z(n347) );
  GTECH_XOR2 U324 ( .A(n326), .B(n353), .Z(n309) );
  GTECH_AND2 U325 ( .A(I_b[6]), .B(I_a[0]), .Z(n353) );
  GTECH_XOR3 U326 ( .A(n354), .B(n355), .C(n323), .Z(n326) );
  GTECH_NAND3 U327 ( .A(I_b[4]), .B(I_a[1]), .C(n356), .Z(n323) );
  GTECH_NOT U328 ( .A(n322), .Z(n355) );
  GTECH_OR_NOT U329 ( .A(n279), .B(I_b[5]), .Z(n322) );
  GTECH_NOT U330 ( .A(n321), .Z(n354) );
  GTECH_OR_NOT U331 ( .A(n242), .B(I_b[4]), .Z(n321) );
  GTECH_XOR3 U332 ( .A(n340), .B(n342), .C(n341), .Z(n336) );
  GTECH_OAI21 U333 ( .A(n357), .B(n358), .C(n359), .Z(n341) );
  GTECH_OAI21 U334 ( .A(n360), .B(n361), .C(n362), .Z(n359) );
  GTECH_NOT U335 ( .A(n361), .Z(n357) );
  GTECH_NOT U336 ( .A(n363), .Z(n342) );
  GTECH_OR_NOT U337 ( .A(n203), .B(I_b[3]), .Z(n363) );
  GTECH_NOT U338 ( .A(n338), .Z(n340) );
  GTECH_OR_NOT U339 ( .A(n180), .B(I_b[2]), .Z(n338) );
  GTECH_NOT U340 ( .A(I_a[4]), .Z(n180) );
  GTECH_NOT U341 ( .A(n364), .Z(n311) );
  GTECH_XOR3 U342 ( .A(n330), .B(n332), .C(n331), .Z(n364) );
  GTECH_OAI21 U343 ( .A(n352), .B(n365), .C(n366), .Z(n331) );
  GTECH_OAI21 U344 ( .A(n350), .B(n367), .C(n351), .Z(n366) );
  GTECH_NOT U345 ( .A(n365), .Z(n350) );
  GTECH_NOT U346 ( .A(n367), .Z(n352) );
  GTECH_NOT U347 ( .A(n368), .Z(n332) );
  GTECH_OR_NOT U348 ( .A(n333), .B(I_a[5]), .Z(n368) );
  GTECH_NOT U349 ( .A(n328), .Z(n330) );
  GTECH_OR_NOT U350 ( .A(n334), .B(I_a[6]), .Z(n328) );
  GTECH_OA22 U351 ( .A(n315), .B(n316), .C(n369), .D(n314), .Z(n344) );
  GTECH_AND_NOT U352 ( .A(n315), .B(n370), .Z(n369) );
  GTECH_XOR3 U353 ( .A(n371), .B(n316), .C(n315), .Z(N145) );
  GTECH_XOR2 U354 ( .A(n372), .B(n356), .Z(n315) );
  GTECH_NOT U355 ( .A(n373), .Z(n356) );
  GTECH_OR_NOT U356 ( .A(n320), .B(I_b[5]), .Z(n373) );
  GTECH_OR_NOT U357 ( .A(n279), .B(I_b[4]), .Z(n372) );
  GTECH_NOT U358 ( .A(n370), .Z(n316) );
  GTECH_XOR2 U359 ( .A(n374), .B(n346), .Z(n370) );
  GTECH_ADD_ABC U360 ( .A(n375), .B(n376), .C(n377), .COUT(n346) );
  GTECH_XOR3 U361 ( .A(n378), .B(n379), .C(n380), .Z(n376) );
  GTECH_OA22 U362 ( .A(n381), .B(n382), .C(n383), .D(n384), .Z(n375) );
  GTECH_AND2 U363 ( .A(n383), .B(n384), .Z(n381) );
  GTECH_XOR4 U364 ( .A(n351), .B(n367), .C(n365), .D(n349), .Z(n374) );
  GTECH_XOR3 U365 ( .A(n360), .B(n362), .C(n361), .Z(n349) );
  GTECH_OAI21 U366 ( .A(n385), .B(n386), .C(n387), .Z(n361) );
  GTECH_NOT U367 ( .A(n388), .Z(n362) );
  GTECH_OR_NOT U368 ( .A(n242), .B(I_b[3]), .Z(n388) );
  GTECH_NOT U369 ( .A(n358), .Z(n360) );
  GTECH_OR_NOT U370 ( .A(n203), .B(I_b[2]), .Z(n358) );
  GTECH_OR_NOT U371 ( .A(n334), .B(I_a[5]), .Z(n365) );
  GTECH_OAI21 U372 ( .A(n380), .B(n389), .C(n390), .Z(n367) );
  GTECH_OAI21 U373 ( .A(n378), .B(n391), .C(n379), .Z(n390) );
  GTECH_NOT U374 ( .A(n391), .Z(n380) );
  GTECH_NOT U375 ( .A(n392), .Z(n351) );
  GTECH_OR_NOT U376 ( .A(n333), .B(I_a[4]), .Z(n392) );
  GTECH_NOT U377 ( .A(n314), .Z(n371) );
  GTECH_NAND3 U378 ( .A(I_a[0]), .B(n393), .C(I_b[4]), .Z(n314) );
  GTECH_XOR2 U379 ( .A(n394), .B(n393), .Z(N144) );
  GTECH_XOR2 U380 ( .A(n395), .B(n396), .Z(n393) );
  GTECH_XOR4 U381 ( .A(n379), .B(n391), .C(n377), .D(n378), .Z(n396) );
  GTECH_NOT U382 ( .A(n389), .Z(n378) );
  GTECH_OR_NOT U383 ( .A(n334), .B(I_a[4]), .Z(n389) );
  GTECH_NOT U384 ( .A(I_b[0]), .Z(n334) );
  GTECH_XOR3 U385 ( .A(n397), .B(n398), .C(n387), .Z(n377) );
  GTECH_NAND3 U386 ( .A(I_b[2]), .B(I_a[1]), .C(n399), .Z(n387) );
  GTECH_NOT U387 ( .A(n386), .Z(n398) );
  GTECH_OR_NOT U388 ( .A(n279), .B(I_b[3]), .Z(n386) );
  GTECH_NOT U389 ( .A(n385), .Z(n397) );
  GTECH_OR_NOT U390 ( .A(n242), .B(I_b[2]), .Z(n385) );
  GTECH_OAI21 U391 ( .A(n400), .B(n401), .C(n402), .Z(n391) );
  GTECH_OAI21 U392 ( .A(n403), .B(n404), .C(n405), .Z(n402) );
  GTECH_NOT U393 ( .A(n404), .Z(n400) );
  GTECH_NOT U394 ( .A(n406), .Z(n379) );
  GTECH_OR_NOT U395 ( .A(n333), .B(I_a[3]), .Z(n406) );
  GTECH_OA22 U396 ( .A(n383), .B(n384), .C(n407), .D(n382), .Z(n395) );
  GTECH_AND_NOT U397 ( .A(n383), .B(n408), .Z(n407) );
  GTECH_AND2 U398 ( .A(I_b[4]), .B(I_a[0]), .Z(n394) );
  GTECH_XOR3 U399 ( .A(n409), .B(n384), .C(n383), .Z(N143) );
  GTECH_XOR2 U400 ( .A(n410), .B(n399), .Z(n383) );
  GTECH_NOT U401 ( .A(n411), .Z(n399) );
  GTECH_OR_NOT U402 ( .A(n320), .B(I_b[3]), .Z(n411) );
  GTECH_NOT U403 ( .A(I_a[0]), .Z(n320) );
  GTECH_OR_NOT U404 ( .A(n279), .B(I_b[2]), .Z(n410) );
  GTECH_NOT U405 ( .A(I_a[1]), .Z(n279) );
  GTECH_NOT U406 ( .A(n408), .Z(n384) );
  GTECH_XOR3 U407 ( .A(n403), .B(n405), .C(n404), .Z(n408) );
  GTECH_OAI21 U408 ( .A(n412), .B(n413), .C(n414), .Z(n404) );
  GTECH_NOT U409 ( .A(n415), .Z(n405) );
  GTECH_OR_NOT U410 ( .A(n242), .B(I_b[1]), .Z(n415) );
  GTECH_NOT U411 ( .A(n401), .Z(n403) );
  GTECH_OR_NOT U412 ( .A(n203), .B(I_b[0]), .Z(n401) );
  GTECH_NOT U413 ( .A(I_a[3]), .Z(n203) );
  GTECH_NOT U414 ( .A(n382), .Z(n409) );
  GTECH_NAND3 U415 ( .A(I_a[0]), .B(n416), .C(I_b[2]), .Z(n382) );
  GTECH_XOR2 U416 ( .A(n417), .B(n416), .Z(N142) );
  GTECH_NOT U417 ( .A(n418), .Z(n416) );
  GTECH_XOR3 U418 ( .A(n419), .B(n420), .C(n414), .Z(n418) );
  GTECH_NAND3 U419 ( .A(n421), .B(I_b[0]), .C(I_a[1]), .Z(n414) );
  GTECH_NOT U420 ( .A(n412), .Z(n420) );
  GTECH_OR_NOT U421 ( .A(n333), .B(I_a[1]), .Z(n412) );
  GTECH_NOT U422 ( .A(n413), .Z(n419) );
  GTECH_OR_NOT U423 ( .A(n242), .B(I_b[0]), .Z(n413) );
  GTECH_NOT U424 ( .A(I_a[2]), .Z(n242) );
  GTECH_AND2 U425 ( .A(I_b[2]), .B(I_a[0]), .Z(n417) );
  GTECH_XOR2 U426 ( .A(n421), .B(n422), .Z(N141) );
  GTECH_AND2 U427 ( .A(I_a[1]), .B(I_b[0]), .Z(n422) );
  GTECH_NOT U428 ( .A(n423), .Z(n421) );
  GTECH_OR_NOT U429 ( .A(n333), .B(I_a[0]), .Z(n423) );
  GTECH_NOT U430 ( .A(I_b[1]), .Z(n333) );
  GTECH_AND2 U431 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

