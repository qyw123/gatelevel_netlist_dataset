
module bcd_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162;

  GTECH_XOR2 U55 ( .A(n87), .B(n88), .Z(sum[9]) );
  GTECH_XOR3 U56 ( .A(b[8]), .B(a[8]), .C(n89), .Z(sum[8]) );
  GTECH_XNOR2 U57 ( .A(n90), .B(n91), .Z(sum[7]) );
  GTECH_AND_NOT U58 ( .A(n92), .B(n93), .Z(n90) );
  GTECH_OAI21 U59 ( .A(n93), .B(n92), .C(n94), .Z(sum[6]) );
  GTECH_OAI21 U60 ( .A(n93), .B(n95), .C(n96), .Z(n94) );
  GTECH_NOT U61 ( .A(n97), .Z(n92) );
  GTECH_XNOR2 U62 ( .A(n95), .B(n93), .Z(sum[5]) );
  GTECH_NOT U63 ( .A(n89), .Z(n93) );
  GTECH_XOR3 U64 ( .A(b[4]), .B(a[4]), .C(n98), .Z(sum[4]) );
  GTECH_XNOR2 U65 ( .A(n99), .B(n100), .Z(sum[3]) );
  GTECH_AND_NOT U66 ( .A(n101), .B(n102), .Z(n99) );
  GTECH_OAI21 U67 ( .A(n102), .B(n101), .C(n103), .Z(sum[2]) );
  GTECH_OAI21 U68 ( .A(n102), .B(n104), .C(n105), .Z(n103) );
  GTECH_NOT U69 ( .A(n106), .Z(n101) );
  GTECH_XNOR2 U70 ( .A(n104), .B(n102), .Z(sum[1]) );
  GTECH_NOT U71 ( .A(n98), .Z(n102) );
  GTECH_XNOR2 U72 ( .A(n107), .B(n108), .Z(sum[15]) );
  GTECH_AND_NOT U73 ( .A(n109), .B(n110), .Z(n107) );
  GTECH_OAI21 U74 ( .A(n110), .B(n109), .C(n111), .Z(sum[14]) );
  GTECH_OAI21 U75 ( .A(n110), .B(n112), .C(n113), .Z(n111) );
  GTECH_NOT U76 ( .A(n114), .Z(n109) );
  GTECH_XNOR2 U77 ( .A(n112), .B(n110), .Z(sum[13]) );
  GTECH_NOT U78 ( .A(cout), .Z(n110) );
  GTECH_XOR3 U79 ( .A(b[12]), .B(a[12]), .C(n115), .Z(sum[12]) );
  GTECH_XNOR2 U80 ( .A(n116), .B(n117), .Z(sum[11]) );
  GTECH_AND_NOT U81 ( .A(n118), .B(n88), .Z(n116) );
  GTECH_OAI21 U82 ( .A(n88), .B(n118), .C(n119), .Z(sum[10]) );
  GTECH_OAI21 U83 ( .A(n88), .B(n120), .C(n121), .Z(n119) );
  GTECH_NOT U84 ( .A(n122), .Z(n118) );
  GTECH_NOT U85 ( .A(n115), .Z(n88) );
  GTECH_XOR3 U86 ( .A(cin), .B(b[0]), .C(a[0]), .Z(sum[0]) );
  GTECH_OAI21 U87 ( .A(n123), .B(n124), .C(n125), .Z(cout) );
  GTECH_OA21 U88 ( .A(n114), .B(n108), .C(n126), .Z(n125) );
  GTECH_OAI21 U89 ( .A(n127), .B(a[15]), .C(b[15]), .Z(n126) );
  GTECH_NOT U90 ( .A(n124), .Z(n127) );
  GTECH_XNOR3 U91 ( .A(b[15]), .B(n123), .C(n124), .Z(n108) );
  GTECH_NOR2 U92 ( .A(n112), .B(n113), .Z(n114) );
  GTECH_XOR3 U93 ( .A(b[14]), .B(a[14]), .C(n128), .Z(n113) );
  GTECH_XOR3 U94 ( .A(b[13]), .B(a[13]), .C(n129), .Z(n112) );
  GTECH_OAI21 U95 ( .A(a[14]), .B(n128), .C(n130), .Z(n124) );
  GTECH_AO21 U96 ( .A(a[14]), .B(n128), .C(b[14]), .Z(n130) );
  GTECH_OA21 U97 ( .A(a[13]), .B(n129), .C(n131), .Z(n128) );
  GTECH_AO21 U98 ( .A(a[13]), .B(n129), .C(b[13]), .Z(n131) );
  GTECH_OA21 U99 ( .A(a[12]), .B(n115), .C(n132), .Z(n129) );
  GTECH_AO21 U100 ( .A(n115), .B(a[12]), .C(b[12]), .Z(n132) );
  GTECH_OAI21 U101 ( .A(n133), .B(n134), .C(n135), .Z(n115) );
  GTECH_OA21 U102 ( .A(n122), .B(n117), .C(n136), .Z(n135) );
  GTECH_OAI21 U103 ( .A(n137), .B(a[11]), .C(b[11]), .Z(n136) );
  GTECH_NOT U104 ( .A(n134), .Z(n137) );
  GTECH_XNOR3 U105 ( .A(b[11]), .B(n133), .C(n134), .Z(n117) );
  GTECH_NOR2 U106 ( .A(n120), .B(n121), .Z(n122) );
  GTECH_XOR3 U107 ( .A(b[10]), .B(a[10]), .C(n138), .Z(n121) );
  GTECH_NOT U108 ( .A(n87), .Z(n120) );
  GTECH_XNOR3 U109 ( .A(b[9]), .B(a[9]), .C(n139), .Z(n87) );
  GTECH_OAI21 U110 ( .A(a[10]), .B(n138), .C(n140), .Z(n134) );
  GTECH_AO21 U111 ( .A(n138), .B(a[10]), .C(b[10]), .Z(n140) );
  GTECH_OA21 U112 ( .A(a[9]), .B(n139), .C(n141), .Z(n138) );
  GTECH_AO21 U113 ( .A(n139), .B(a[9]), .C(b[9]), .Z(n141) );
  GTECH_OA21 U114 ( .A(a[8]), .B(n89), .C(n142), .Z(n139) );
  GTECH_AO21 U115 ( .A(n89), .B(a[8]), .C(b[8]), .Z(n142) );
  GTECH_OAI21 U116 ( .A(n143), .B(n144), .C(n145), .Z(n89) );
  GTECH_OA21 U117 ( .A(n97), .B(n91), .C(n146), .Z(n145) );
  GTECH_OAI21 U118 ( .A(n147), .B(a[7]), .C(b[7]), .Z(n146) );
  GTECH_NOT U119 ( .A(n144), .Z(n147) );
  GTECH_XNOR3 U120 ( .A(b[7]), .B(n143), .C(n144), .Z(n91) );
  GTECH_NOR2 U121 ( .A(n95), .B(n96), .Z(n97) );
  GTECH_XOR3 U122 ( .A(b[6]), .B(a[6]), .C(n148), .Z(n96) );
  GTECH_XOR3 U123 ( .A(b[5]), .B(a[5]), .C(n149), .Z(n95) );
  GTECH_OAI21 U124 ( .A(a[6]), .B(n148), .C(n150), .Z(n144) );
  GTECH_AO21 U125 ( .A(n148), .B(a[6]), .C(b[6]), .Z(n150) );
  GTECH_OA21 U126 ( .A(a[5]), .B(n149), .C(n151), .Z(n148) );
  GTECH_AO21 U127 ( .A(n149), .B(a[5]), .C(b[5]), .Z(n151) );
  GTECH_OA21 U128 ( .A(a[4]), .B(n98), .C(n152), .Z(n149) );
  GTECH_AO21 U129 ( .A(n98), .B(a[4]), .C(b[4]), .Z(n152) );
  GTECH_OAI21 U130 ( .A(n153), .B(n154), .C(n155), .Z(n98) );
  GTECH_OA21 U131 ( .A(n106), .B(n100), .C(n156), .Z(n155) );
  GTECH_OAI21 U132 ( .A(n157), .B(a[3]), .C(b[3]), .Z(n156) );
  GTECH_NOT U133 ( .A(n154), .Z(n157) );
  GTECH_XNOR3 U134 ( .A(b[3]), .B(n153), .C(n154), .Z(n100) );
  GTECH_NOR2 U135 ( .A(n104), .B(n105), .Z(n106) );
  GTECH_XOR3 U136 ( .A(b[2]), .B(a[2]), .C(n158), .Z(n105) );
  GTECH_XOR3 U137 ( .A(b[1]), .B(a[1]), .C(n159), .Z(n104) );
  GTECH_OAI21 U138 ( .A(a[2]), .B(n158), .C(n160), .Z(n154) );
  GTECH_AO21 U139 ( .A(n158), .B(a[2]), .C(b[2]), .Z(n160) );
  GTECH_OA21 U140 ( .A(a[1]), .B(n159), .C(n161), .Z(n158) );
  GTECH_AO21 U141 ( .A(n159), .B(a[1]), .C(b[1]), .Z(n161) );
  GTECH_OA21 U142 ( .A(b[0]), .B(a[0]), .C(n162), .Z(n159) );
  GTECH_AO21 U143 ( .A(a[0]), .B(b[0]), .C(cin), .Z(n162) );
  GTECH_NOT U144 ( .A(a[3]), .Z(n153) );
  GTECH_NOT U145 ( .A(a[7]), .Z(n143) );
  GTECH_NOT U146 ( .A(a[11]), .Z(n133) );
  GTECH_NOT U147 ( .A(a[15]), .Z(n123) );
endmodule

