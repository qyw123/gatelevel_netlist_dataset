
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n128, n129, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK2S Cntr_reg_0_ ( .J(n129), .K(n129), .TI(N14), .TE(N18), .CP(clk), 
        .CD(n128), .Q(Cntr[0]), .QN(n353) );
  GTECH_FJK2S Cntr_reg_1_ ( .J(n129), .K(n129), .TI(N15), .TE(N18), .CP(clk), 
        .CD(n128), .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK2S Cntr_reg_2_ ( .J(n129), .K(n129), .TI(N16), .TE(N18), .CP(clk), 
        .CD(n128), .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK2S Cntr_reg_3_ ( .J(n129), .K(n129), .TI(N17), .TE(N18), .CP(clk), 
        .CD(n128), .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK2S Cntr_reg_4_ ( .J(n129), .K(n129), .TI(N19), .TE(N18), .CP(clk), 
        .CD(n128), .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK2S A_reg_16_ ( .J(n129), .K(n129), .TI(N42), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[16]), .QN(n370) );
  GTECH_FJK2S A_reg_15_ ( .J(n129), .K(n129), .TI(N42), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[15]), .QN(n369) );
  GTECH_FJK2S A_reg_14_ ( .J(n129), .K(n129), .TI(N39), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[14]), .QN(n368) );
  GTECH_FJK2S A_reg_13_ ( .J(n129), .K(n129), .TI(N38), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[13]), .QN(n367) );
  GTECH_FJK2S A_reg_12_ ( .J(n129), .K(n129), .TI(N37), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[12]), .QN(n366) );
  GTECH_FJK2S A_reg_11_ ( .J(n129), .K(n129), .TI(N36), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[11]), .QN(n365) );
  GTECH_FJK2S A_reg_10_ ( .J(n129), .K(n129), .TI(N35), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[10]), .QN(n364) );
  GTECH_FJK2S A_reg_9_ ( .J(n129), .K(n129), .TI(N34), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[9]), .QN(n363) );
  GTECH_FJK2S A_reg_8_ ( .J(n129), .K(n129), .TI(N33), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[8]), .QN(n362) );
  GTECH_FJK2S A_reg_7_ ( .J(n129), .K(n129), .TI(N32), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[7]), .QN(n361) );
  GTECH_FJK2S A_reg_6_ ( .J(n129), .K(n129), .TI(N31), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[6]), .QN(n360) );
  GTECH_FJK2S A_reg_5_ ( .J(n129), .K(n129), .TI(N30), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[5]), .QN(n359) );
  GTECH_FJK2S A_reg_4_ ( .J(n129), .K(n129), .TI(N29), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[4]), .QN(n358) );
  GTECH_FJK2S A_reg_3_ ( .J(n129), .K(n129), .TI(N28), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[3]), .QN(n357) );
  GTECH_FJK2S A_reg_2_ ( .J(n129), .K(n129), .TI(N27), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[2]), .QN(n356) );
  GTECH_FJK2S A_reg_1_ ( .J(n129), .K(n129), .TI(N26), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[1]), .QN(n355) );
  GTECH_FJK2S A_reg_0_ ( .J(n129), .K(n129), .TI(N25), .TE(N41), .CP(clk), 
        .CD(n128), .Q(A[0]), .QN(n354) );
  GTECH_FJK2S Prod_reg_0_ ( .J(n129), .K(n129), .TI(N82), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[0]), .QN(n10) );
  GTECH_FJK2S Prod_reg_18_ ( .J(n129), .K(n129), .TI(N100), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK2S Prod_reg_17_ ( .J(n129), .K(n129), .TI(N99), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[17]), .QN(n12) );
  GTECH_FJK2S Prod_reg_16_ ( .J(n129), .K(n129), .TI(N98), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[16]), .QN(n13) );
  GTECH_FJK2S Prod_reg_15_ ( .J(n129), .K(n129), .TI(N97), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[15]), .QN(n14) );
  GTECH_FJK2S Prod_reg_14_ ( .J(n129), .K(n129), .TI(N96), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[14]), .QN(n15) );
  GTECH_FJK2S Prod_reg_13_ ( .J(n129), .K(n129), .TI(N95), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[13]), .QN(n16) );
  GTECH_FJK2S Prod_reg_12_ ( .J(n129), .K(n129), .TI(N94), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[12]), .QN(n17) );
  GTECH_FJK2S Prod_reg_11_ ( .J(n129), .K(n129), .TI(N93), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[11]), .QN(n18) );
  GTECH_FJK2S Prod_reg_10_ ( .J(n129), .K(n129), .TI(N92), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[10]), .QN(n19) );
  GTECH_FJK2S Prod_reg_9_ ( .J(n129), .K(n129), .TI(N91), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[9]), .QN(n20) );
  GTECH_FJK2S Prod_reg_8_ ( .J(n129), .K(n129), .TI(N90), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[8]), .QN(n21) );
  GTECH_FJK2S Prod_reg_7_ ( .J(n129), .K(n129), .TI(N89), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[7]), .QN(n22) );
  GTECH_FJK2S Prod_reg_6_ ( .J(n129), .K(n129), .TI(N88), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[6]), .QN(n23) );
  GTECH_FJK2S Prod_reg_5_ ( .J(n129), .K(n129), .TI(N87), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[5]), .QN(n24) );
  GTECH_FJK2S Prod_reg_4_ ( .J(n129), .K(n129), .TI(N86), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[4]), .QN(n25) );
  GTECH_FJK2S Prod_reg_3_ ( .J(n129), .K(n129), .TI(N85), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[3]), .QN(n26) );
  GTECH_FJK2S Prod_reg_2_ ( .J(n129), .K(n129), .TI(N84), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[2]), .QN(n27) );
  GTECH_FJK2S Prod_reg_1_ ( .J(n129), .K(n129), .TI(N83), .TE(N115), .CP(clk), 
        .CD(n128), .Q(Prod[1]), .QN(n28) );
  GTECH_FJK2S Prod_reg_19_ ( .J(n129), .K(n129), .TI(N101), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK2S Prod_reg_33_ ( .J(n129), .K(n129), .TI(N116), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK2S Prod_reg_32_ ( .J(n129), .K(n129), .TI(N116), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK2S Prod_reg_31_ ( .J(n129), .K(n129), .TI(N113), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK2S Prod_reg_30_ ( .J(n129), .K(n129), .TI(N112), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK2S Prod_reg_29_ ( .J(n129), .K(n129), .TI(N111), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK2S Prod_reg_28_ ( .J(n129), .K(n129), .TI(N110), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK2S Prod_reg_27_ ( .J(n129), .K(n129), .TI(N109), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK2S Prod_reg_26_ ( .J(n129), .K(n129), .TI(N108), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK2S Prod_reg_25_ ( .J(n129), .K(n129), .TI(N107), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK2S Prod_reg_24_ ( .J(n129), .K(n129), .TI(N106), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK2S Prod_reg_23_ ( .J(n129), .K(n129), .TI(N105), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK2S Prod_reg_22_ ( .J(n129), .K(n129), .TI(N104), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK2S Prod_reg_21_ ( .J(n129), .K(n129), .TI(N103), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK2S Prod_reg_20_ ( .J(n129), .K(n129), .TI(N102), .TE(N115), .CP(clk), .CD(n128), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK2S P_reg_31_ ( .J(n129), .K(n129), .TI(N152), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[31]) );
  GTECH_FJK2S P_reg_30_ ( .J(n129), .K(n129), .TI(N150), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[30]) );
  GTECH_FJK2S P_reg_29_ ( .J(n129), .K(n129), .TI(N149), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[29]) );
  GTECH_FJK2S P_reg_28_ ( .J(n129), .K(n129), .TI(N148), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[28]) );
  GTECH_FJK2S P_reg_27_ ( .J(n129), .K(n129), .TI(N147), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[27]) );
  GTECH_FJK2S P_reg_26_ ( .J(n129), .K(n129), .TI(N146), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[26]) );
  GTECH_FJK2S P_reg_25_ ( .J(n129), .K(n129), .TI(N145), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[25]) );
  GTECH_FJK2S P_reg_24_ ( .J(n129), .K(n129), .TI(N144), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[24]) );
  GTECH_FJK2S P_reg_23_ ( .J(n129), .K(n129), .TI(N143), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[23]) );
  GTECH_FJK2S P_reg_22_ ( .J(n129), .K(n129), .TI(N142), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[22]) );
  GTECH_FJK2S P_reg_21_ ( .J(n129), .K(n129), .TI(N141), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[21]) );
  GTECH_FJK2S P_reg_20_ ( .J(n129), .K(n129), .TI(N140), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[20]) );
  GTECH_FJK2S P_reg_19_ ( .J(n129), .K(n129), .TI(N139), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[19]) );
  GTECH_FJK2S P_reg_18_ ( .J(n129), .K(n129), .TI(N138), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[18]) );
  GTECH_FJK2S P_reg_17_ ( .J(n129), .K(n129), .TI(N137), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[17]) );
  GTECH_FJK2S P_reg_16_ ( .J(n129), .K(n129), .TI(N136), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[16]) );
  GTECH_FJK2S P_reg_15_ ( .J(n129), .K(n129), .TI(N135), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[15]) );
  GTECH_FJK2S P_reg_14_ ( .J(n129), .K(n129), .TI(N134), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[14]) );
  GTECH_FJK2S P_reg_13_ ( .J(n129), .K(n129), .TI(N133), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[13]) );
  GTECH_FJK2S P_reg_12_ ( .J(n129), .K(n129), .TI(N132), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[12]) );
  GTECH_FJK2S P_reg_11_ ( .J(n129), .K(n129), .TI(N131), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[11]) );
  GTECH_FJK2S P_reg_10_ ( .J(n129), .K(n129), .TI(N130), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[10]) );
  GTECH_FJK2S P_reg_9_ ( .J(n129), .K(n129), .TI(N129), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[9]) );
  GTECH_FJK2S P_reg_8_ ( .J(n129), .K(n129), .TI(N128), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[8]) );
  GTECH_FJK2S P_reg_7_ ( .J(n129), .K(n129), .TI(N127), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[7]) );
  GTECH_FJK2S P_reg_6_ ( .J(n129), .K(n129), .TI(N126), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[6]) );
  GTECH_FJK2S P_reg_5_ ( .J(n129), .K(n129), .TI(N125), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[5]) );
  GTECH_FJK2S P_reg_4_ ( .J(n129), .K(n129), .TI(N124), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[4]) );
  GTECH_FJK2S P_reg_3_ ( .J(n129), .K(n129), .TI(N123), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[3]) );
  GTECH_FJK2S P_reg_2_ ( .J(n129), .K(n129), .TI(N122), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[2]) );
  GTECH_FJK2S P_reg_1_ ( .J(n129), .K(n129), .TI(N121), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[1]) );
  GTECH_FJK2S P_reg_0_ ( .J(n129), .K(n129), .TI(N120), .TE(N151), .CP(clk), 
        .CD(n128), .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U355 ( .Z(n129) );
  GTECH_ONE U356 ( .Z(n128) );
  GTECH_NOT U357 ( .A(n371), .Z(N99) );
  GTECH_AOI222 U358 ( .A(n372), .B(n373), .C(n374), .D(n375), .E(n376), .F(
        n377), .Z(n371) );
  GTECH_NOT U359 ( .A(n378), .Z(N98) );
  GTECH_AOI222 U360 ( .A(n374), .B(n379), .C(n380), .D(n381), .E(R[15]), .F(
        n382), .Z(n378) );
  GTECH_NAND2 U361 ( .A(n383), .B(n384), .Z(n380) );
  GTECH_AO22 U362 ( .A(n385), .B(n386), .C(R[14]), .D(n382), .Z(N97) );
  GTECH_AO22 U363 ( .A(n385), .B(n387), .C(R[13]), .D(n382), .Z(N96) );
  GTECH_AO22 U364 ( .A(n385), .B(n388), .C(R[12]), .D(n382), .Z(N95) );
  GTECH_AO22 U365 ( .A(n385), .B(n389), .C(R[11]), .D(n382), .Z(N94) );
  GTECH_AO22 U366 ( .A(n385), .B(n390), .C(R[10]), .D(n382), .Z(N93) );
  GTECH_AO22 U367 ( .A(n385), .B(n391), .C(R[9]), .D(n382), .Z(N92) );
  GTECH_AO22 U368 ( .A(n385), .B(n392), .C(R[8]), .D(n382), .Z(N91) );
  GTECH_AO22 U369 ( .A(n385), .B(n393), .C(R[7]), .D(n382), .Z(N90) );
  GTECH_AO22 U370 ( .A(n385), .B(n394), .C(R[6]), .D(n382), .Z(N89) );
  GTECH_AO22 U371 ( .A(n385), .B(n395), .C(R[5]), .D(n382), .Z(N88) );
  GTECH_AO22 U372 ( .A(n385), .B(n396), .C(R[4]), .D(n382), .Z(N87) );
  GTECH_AO22 U373 ( .A(n385), .B(n397), .C(R[3]), .D(n382), .Z(N86) );
  GTECH_AO22 U374 ( .A(n385), .B(n398), .C(R[2]), .D(n382), .Z(N85) );
  GTECH_AO22 U375 ( .A(n385), .B(n399), .C(R[1]), .D(n382), .Z(N84) );
  GTECH_AO22 U376 ( .A(n385), .B(n400), .C(R[0]), .D(n382), .Z(N83) );
  GTECH_AND2 U377 ( .A(M[15]), .B(n382), .Z(N42) );
  GTECH_AND2 U378 ( .A(M[14]), .B(n382), .Z(N39) );
  GTECH_AND2 U379 ( .A(M[13]), .B(n382), .Z(N38) );
  GTECH_AND2 U380 ( .A(M[12]), .B(n382), .Z(N37) );
  GTECH_AND2 U381 ( .A(M[11]), .B(n382), .Z(N36) );
  GTECH_AND2 U382 ( .A(M[10]), .B(n382), .Z(N35) );
  GTECH_AND2 U383 ( .A(M[9]), .B(n382), .Z(N34) );
  GTECH_AND2 U384 ( .A(M[8]), .B(n382), .Z(N33) );
  GTECH_AND2 U385 ( .A(M[7]), .B(n382), .Z(N32) );
  GTECH_AND2 U386 ( .A(M[6]), .B(n382), .Z(N31) );
  GTECH_AND2 U387 ( .A(M[5]), .B(n382), .Z(N30) );
  GTECH_AND2 U388 ( .A(M[4]), .B(n382), .Z(N29) );
  GTECH_AND2 U389 ( .A(M[3]), .B(n382), .Z(N28) );
  GTECH_AND2 U390 ( .A(M[2]), .B(n382), .Z(N27) );
  GTECH_AND2 U391 ( .A(M[1]), .B(n382), .Z(N26) );
  GTECH_AND2 U392 ( .A(M[0]), .B(n382), .Z(N25) );
  GTECH_NOT U393 ( .A(n401), .Z(n382) );
  GTECH_NAND2 U394 ( .A(n401), .B(n402), .Z(N19) );
  GTECH_NAND3 U395 ( .A(n403), .B(n404), .C(n385), .Z(n402) );
  GTECH_NAND3 U396 ( .A(n405), .B(n406), .C(n407), .Z(N18) );
  GTECH_AND2 U397 ( .A(n385), .B(n408), .Z(N17) );
  GTECH_OAI21 U398 ( .A(n8), .B(n409), .C(n403), .Z(n408) );
  GTECH_AND2 U399 ( .A(n385), .B(n410), .Z(N16) );
  GTECH_OAI21 U400 ( .A(n7), .B(n411), .C(n412), .Z(n410) );
  GTECH_NOT U401 ( .A(n413), .Z(N152) );
  GTECH_AOI222 U402 ( .A(n414), .B(n415), .C(n416), .D(n417), .E(n418), .F(
        n419), .Z(n413) );
  GTECH_NAND2 U403 ( .A(n406), .B(n420), .Z(N151) );
  GTECH_NOT U404 ( .A(n421), .Z(N150) );
  GTECH_AOI222 U405 ( .A(n422), .B(n414), .C(n416), .D(n423), .E(n418), .F(
        n424), .Z(n421) );
  GTECH_MUX2 U406 ( .A(n425), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND2 U407 ( .A(n385), .B(n426), .Z(n425) );
  GTECH_NOT U408 ( .A(n427), .Z(N149) );
  GTECH_AOI222 U409 ( .A(n428), .B(n414), .C(n416), .D(n429), .E(n418), .F(
        n430), .Z(n427) );
  GTECH_NOT U410 ( .A(n431), .Z(N148) );
  GTECH_AOI222 U411 ( .A(n432), .B(n414), .C(n416), .D(n433), .E(n418), .F(
        n434), .Z(n431) );
  GTECH_NOT U412 ( .A(n435), .Z(N147) );
  GTECH_AOI222 U413 ( .A(n436), .B(n414), .C(n416), .D(n437), .E(n418), .F(
        n438), .Z(n435) );
  GTECH_NOT U414 ( .A(n439), .Z(N146) );
  GTECH_AOI222 U415 ( .A(n440), .B(n414), .C(n416), .D(n441), .E(n418), .F(
        n442), .Z(n439) );
  GTECH_NOT U416 ( .A(n443), .Z(N145) );
  GTECH_AOI222 U417 ( .A(n444), .B(n414), .C(n416), .D(n445), .E(n418), .F(
        n446), .Z(n443) );
  GTECH_NOT U418 ( .A(n447), .Z(N144) );
  GTECH_AOI222 U419 ( .A(n448), .B(n414), .C(n416), .D(n449), .E(n418), .F(
        n450), .Z(n447) );
  GTECH_NOT U420 ( .A(n451), .Z(N143) );
  GTECH_AOI222 U421 ( .A(n452), .B(n414), .C(n416), .D(n453), .E(n418), .F(
        n454), .Z(n451) );
  GTECH_NOT U422 ( .A(n455), .Z(N142) );
  GTECH_AOI222 U423 ( .A(n456), .B(n414), .C(n416), .D(n457), .E(n418), .F(
        n458), .Z(n455) );
  GTECH_NOT U424 ( .A(n459), .Z(N141) );
  GTECH_AOI222 U425 ( .A(n460), .B(n414), .C(n416), .D(n461), .E(n418), .F(
        n462), .Z(n459) );
  GTECH_NOT U426 ( .A(n463), .Z(N140) );
  GTECH_AOI222 U427 ( .A(n464), .B(n414), .C(n416), .D(n465), .E(n418), .F(
        n466), .Z(n463) );
  GTECH_NOT U428 ( .A(n467), .Z(N14) );
  GTECH_NAND2 U429 ( .A(n385), .B(n353), .Z(n467) );
  GTECH_NOT U430 ( .A(n468), .Z(N139) );
  GTECH_AOI222 U431 ( .A(n469), .B(n414), .C(n416), .D(n470), .E(n418), .F(
        n471), .Z(n468) );
  GTECH_NOT U432 ( .A(n472), .Z(N138) );
  GTECH_AOI222 U433 ( .A(n473), .B(n414), .C(n416), .D(n474), .E(n418), .F(
        n475), .Z(n472) );
  GTECH_NOT U434 ( .A(n476), .Z(N137) );
  GTECH_AOI222 U435 ( .A(n477), .B(n414), .C(n416), .D(n478), .E(n418), .F(
        n479), .Z(n476) );
  GTECH_NOT U436 ( .A(n480), .Z(N136) );
  GTECH_AOI222 U437 ( .A(n414), .B(n373), .C(n416), .D(n375), .E(n418), .F(
        n377), .Z(n480) );
  GTECH_NOT U438 ( .A(n481), .Z(n377) );
  GTECH_XOR2 U439 ( .A(n482), .B(n483), .Z(n481) );
  GTECH_NOT U440 ( .A(n484), .Z(n483) );
  GTECH_NOT U441 ( .A(n485), .Z(n416) );
  GTECH_NOT U442 ( .A(n486), .Z(n373) );
  GTECH_XOR2 U443 ( .A(n482), .B(n487), .Z(n486) );
  GTECH_NOT U444 ( .A(n488), .Z(n487) );
  GTECH_XOR2 U445 ( .A(n375), .B(n355), .Z(n482) );
  GTECH_OAI21 U446 ( .A(n12), .B(n485), .C(n489), .Z(N135) );
  GTECH_OAI21 U447 ( .A(n418), .B(n414), .C(n381), .Z(n489) );
  GTECH_OAI21 U448 ( .A(n12), .B(n490), .C(n484), .Z(n381) );
  GTECH_NOT U449 ( .A(n491), .Z(n414) );
  GTECH_NAND3 U450 ( .A(n28), .B(n492), .C(N155), .Z(n491) );
  GTECH_NOT U451 ( .A(n493), .Z(n418) );
  GTECH_NAND3 U452 ( .A(n10), .B(n494), .C(N155), .Z(n493) );
  GTECH_NAND2 U453 ( .A(n495), .B(N155), .Z(n485) );
  GTECH_XOR2 U454 ( .A(n492), .B(n28), .Z(n495) );
  GTECH_AND2 U455 ( .A(N155), .B(n386), .Z(N134) );
  GTECH_NOT U456 ( .A(n13), .Z(n386) );
  GTECH_AND2 U457 ( .A(N155), .B(n387), .Z(N133) );
  GTECH_NOT U458 ( .A(n14), .Z(n387) );
  GTECH_AND2 U459 ( .A(N155), .B(n388), .Z(N132) );
  GTECH_NOT U460 ( .A(n15), .Z(n388) );
  GTECH_AND2 U461 ( .A(N155), .B(n389), .Z(N131) );
  GTECH_NOT U462 ( .A(n16), .Z(n389) );
  GTECH_AND2 U463 ( .A(N155), .B(n390), .Z(N130) );
  GTECH_NOT U464 ( .A(n17), .Z(n390) );
  GTECH_AND2 U465 ( .A(N155), .B(n391), .Z(N129) );
  GTECH_NOT U466 ( .A(n18), .Z(n391) );
  GTECH_AND2 U467 ( .A(N155), .B(n392), .Z(N128) );
  GTECH_NOT U468 ( .A(n19), .Z(n392) );
  GTECH_AND2 U469 ( .A(N155), .B(n393), .Z(N127) );
  GTECH_NOT U470 ( .A(n20), .Z(n393) );
  GTECH_AND2 U471 ( .A(N155), .B(n394), .Z(N126) );
  GTECH_NOT U472 ( .A(n21), .Z(n394) );
  GTECH_AND2 U473 ( .A(N155), .B(n395), .Z(N125) );
  GTECH_NOT U474 ( .A(n22), .Z(n395) );
  GTECH_AND2 U475 ( .A(N155), .B(n396), .Z(N124) );
  GTECH_NOT U476 ( .A(n23), .Z(n396) );
  GTECH_AND2 U477 ( .A(N155), .B(n397), .Z(N123) );
  GTECH_NOT U478 ( .A(n24), .Z(n397) );
  GTECH_AND2 U479 ( .A(N155), .B(n398), .Z(N122) );
  GTECH_NOT U480 ( .A(n25), .Z(n398) );
  GTECH_AND2 U481 ( .A(N155), .B(n399), .Z(N121) );
  GTECH_NOT U482 ( .A(n26), .Z(n399) );
  GTECH_AND2 U483 ( .A(N155), .B(n400), .Z(N120) );
  GTECH_NOT U484 ( .A(n27), .Z(n400) );
  GTECH_NOT U485 ( .A(n420), .Z(N155) );
  GTECH_NAND4 U486 ( .A(n8), .B(n7), .C(n9), .D(n496), .Z(n420) );
  GTECH_AND3 U487 ( .A(n406), .B(n426), .C(n6), .Z(n496) );
  GTECH_NOT U488 ( .A(n353), .Z(n426) );
  GTECH_NOT U489 ( .A(n497), .Z(N116) );
  GTECH_AOI222 U490 ( .A(n374), .B(n417), .C(n376), .D(n419), .E(n415), .F(
        n372), .Z(n497) );
  GTECH_XOR2 U491 ( .A(n498), .B(n499), .Z(n415) );
  GTECH_ADD_ABC U492 ( .A(n369), .B(n31), .C(n500), .COUT(n499) );
  GTECH_XOR2 U493 ( .A(n501), .B(n498), .Z(n419) );
  GTECH_XOR2 U494 ( .A(n417), .B(n370), .Z(n498) );
  GTECH_NAND2 U495 ( .A(n502), .B(n503), .Z(n501) );
  GTECH_OAI21 U496 ( .A(n369), .B(n423), .C(n504), .Z(n503) );
  GTECH_OR_NOT U497 ( .A(n31), .B(n369), .Z(n502) );
  GTECH_NOT U498 ( .A(n30), .Z(n417) );
  GTECH_NAND2 U499 ( .A(n407), .B(n505), .Z(N115) );
  GTECH_NOT U500 ( .A(N41), .Z(n505) );
  GTECH_NAND2 U501 ( .A(n406), .B(n401), .Z(N41) );
  GTECH_NAND2 U502 ( .A(Ld), .B(n406), .Z(n401) );
  GTECH_NOT U503 ( .A(n506), .Z(N113) );
  GTECH_AOI222 U504 ( .A(n374), .B(n423), .C(n376), .D(n424), .E(n422), .F(
        n372), .Z(n506) );
  GTECH_XOR2 U505 ( .A(n507), .B(n500), .Z(n422) );
  GTECH_ADD_ABC U506 ( .A(n368), .B(n32), .C(n508), .COUT(n500) );
  GTECH_NOT U507 ( .A(n509), .Z(n424) );
  GTECH_XOR2 U508 ( .A(n507), .B(n510), .Z(n509) );
  GTECH_NOT U509 ( .A(n504), .Z(n510) );
  GTECH_OAI21 U510 ( .A(n32), .B(n511), .C(n512), .Z(n504) );
  GTECH_OAI21 U511 ( .A(n368), .B(n429), .C(n513), .Z(n512) );
  GTECH_NOT U512 ( .A(n368), .Z(n511) );
  GTECH_XOR2 U513 ( .A(n423), .B(n369), .Z(n507) );
  GTECH_NOT U514 ( .A(n31), .Z(n423) );
  GTECH_NOT U515 ( .A(n514), .Z(N112) );
  GTECH_AOI222 U516 ( .A(n374), .B(n429), .C(n376), .D(n430), .E(n428), .F(
        n372), .Z(n514) );
  GTECH_XOR2 U517 ( .A(n515), .B(n508), .Z(n428) );
  GTECH_ADD_ABC U518 ( .A(n367), .B(n33), .C(n516), .COUT(n508) );
  GTECH_NOT U519 ( .A(n517), .Z(n430) );
  GTECH_XOR2 U520 ( .A(n515), .B(n518), .Z(n517) );
  GTECH_NOT U521 ( .A(n513), .Z(n518) );
  GTECH_OAI21 U522 ( .A(n33), .B(n519), .C(n520), .Z(n513) );
  GTECH_OAI21 U523 ( .A(n367), .B(n433), .C(n521), .Z(n520) );
  GTECH_NOT U524 ( .A(n367), .Z(n519) );
  GTECH_XOR2 U525 ( .A(n429), .B(n368), .Z(n515) );
  GTECH_NOT U526 ( .A(n32), .Z(n429) );
  GTECH_NOT U527 ( .A(n522), .Z(N111) );
  GTECH_AOI222 U528 ( .A(n374), .B(n433), .C(n376), .D(n434), .E(n432), .F(
        n372), .Z(n522) );
  GTECH_XOR2 U529 ( .A(n523), .B(n516), .Z(n432) );
  GTECH_ADD_ABC U530 ( .A(n34), .B(n366), .C(n524), .COUT(n516) );
  GTECH_NOT U531 ( .A(n525), .Z(n434) );
  GTECH_XOR2 U532 ( .A(n523), .B(n526), .Z(n525) );
  GTECH_NOT U533 ( .A(n521), .Z(n526) );
  GTECH_OAI21 U534 ( .A(n34), .B(n527), .C(n528), .Z(n521) );
  GTECH_OAI21 U535 ( .A(n366), .B(n437), .C(n529), .Z(n528) );
  GTECH_XOR2 U536 ( .A(n433), .B(n367), .Z(n523) );
  GTECH_NOT U537 ( .A(n33), .Z(n433) );
  GTECH_NOT U538 ( .A(n530), .Z(N110) );
  GTECH_AOI222 U539 ( .A(n374), .B(n437), .C(n376), .D(n438), .E(n436), .F(
        n372), .Z(n530) );
  GTECH_XOR2 U540 ( .A(n531), .B(n524), .Z(n436) );
  GTECH_ADD_ABC U541 ( .A(n35), .B(n365), .C(n532), .COUT(n524) );
  GTECH_NOT U542 ( .A(n533), .Z(n438) );
  GTECH_XOR2 U543 ( .A(n531), .B(n534), .Z(n533) );
  GTECH_NOT U544 ( .A(n529), .Z(n534) );
  GTECH_OAI21 U545 ( .A(n35), .B(n535), .C(n536), .Z(n529) );
  GTECH_OAI21 U546 ( .A(n365), .B(n441), .C(n537), .Z(n536) );
  GTECH_XOR2 U547 ( .A(n527), .B(n34), .Z(n531) );
  GTECH_NOT U548 ( .A(n366), .Z(n527) );
  GTECH_NOT U549 ( .A(n34), .Z(n437) );
  GTECH_NOT U550 ( .A(n538), .Z(N109) );
  GTECH_AOI222 U551 ( .A(n374), .B(n441), .C(n376), .D(n442), .E(n440), .F(
        n372), .Z(n538) );
  GTECH_XOR2 U552 ( .A(n539), .B(n532), .Z(n440) );
  GTECH_ADD_ABC U553 ( .A(n36), .B(n364), .C(n540), .COUT(n532) );
  GTECH_NOT U554 ( .A(n541), .Z(n442) );
  GTECH_XOR2 U555 ( .A(n539), .B(n542), .Z(n541) );
  GTECH_NOT U556 ( .A(n537), .Z(n542) );
  GTECH_OAI21 U557 ( .A(n36), .B(n543), .C(n544), .Z(n537) );
  GTECH_OAI21 U558 ( .A(n364), .B(n445), .C(n545), .Z(n544) );
  GTECH_XOR2 U559 ( .A(n535), .B(n35), .Z(n539) );
  GTECH_NOT U560 ( .A(n365), .Z(n535) );
  GTECH_NOT U561 ( .A(n35), .Z(n441) );
  GTECH_NOT U562 ( .A(n546), .Z(N108) );
  GTECH_AOI222 U563 ( .A(n374), .B(n445), .C(n376), .D(n446), .E(n444), .F(
        n372), .Z(n546) );
  GTECH_XOR2 U564 ( .A(n547), .B(n540), .Z(n444) );
  GTECH_ADD_ABC U565 ( .A(n37), .B(n363), .C(n548), .COUT(n540) );
  GTECH_NOT U566 ( .A(n549), .Z(n446) );
  GTECH_XOR2 U567 ( .A(n547), .B(n550), .Z(n549) );
  GTECH_NOT U568 ( .A(n545), .Z(n550) );
  GTECH_OAI21 U569 ( .A(n37), .B(n551), .C(n552), .Z(n545) );
  GTECH_OAI21 U570 ( .A(n363), .B(n449), .C(n553), .Z(n552) );
  GTECH_XOR2 U571 ( .A(n543), .B(n36), .Z(n547) );
  GTECH_NOT U572 ( .A(n364), .Z(n543) );
  GTECH_NOT U573 ( .A(n36), .Z(n445) );
  GTECH_NOT U574 ( .A(n554), .Z(N107) );
  GTECH_AOI222 U575 ( .A(n374), .B(n449), .C(n376), .D(n450), .E(n448), .F(
        n372), .Z(n554) );
  GTECH_XOR2 U576 ( .A(n555), .B(n548), .Z(n448) );
  GTECH_ADD_ABC U577 ( .A(n38), .B(n362), .C(n556), .COUT(n548) );
  GTECH_NOT U578 ( .A(n557), .Z(n450) );
  GTECH_XOR2 U579 ( .A(n555), .B(n558), .Z(n557) );
  GTECH_NOT U580 ( .A(n553), .Z(n558) );
  GTECH_OAI21 U581 ( .A(n38), .B(n559), .C(n560), .Z(n553) );
  GTECH_OAI21 U582 ( .A(n362), .B(n453), .C(n561), .Z(n560) );
  GTECH_XOR2 U583 ( .A(n551), .B(n37), .Z(n555) );
  GTECH_NOT U584 ( .A(n363), .Z(n551) );
  GTECH_NOT U585 ( .A(n37), .Z(n449) );
  GTECH_NOT U586 ( .A(n562), .Z(N106) );
  GTECH_AOI222 U587 ( .A(n374), .B(n453), .C(n376), .D(n454), .E(n452), .F(
        n372), .Z(n562) );
  GTECH_XOR2 U588 ( .A(n563), .B(n556), .Z(n452) );
  GTECH_ADD_ABC U589 ( .A(n39), .B(n361), .C(n564), .COUT(n556) );
  GTECH_NOT U590 ( .A(n565), .Z(n454) );
  GTECH_XOR2 U591 ( .A(n563), .B(n566), .Z(n565) );
  GTECH_NOT U592 ( .A(n561), .Z(n566) );
  GTECH_OAI21 U593 ( .A(n39), .B(n567), .C(n568), .Z(n561) );
  GTECH_OAI21 U594 ( .A(n361), .B(n457), .C(n569), .Z(n568) );
  GTECH_XOR2 U595 ( .A(n559), .B(n38), .Z(n563) );
  GTECH_NOT U596 ( .A(n362), .Z(n559) );
  GTECH_NOT U597 ( .A(n38), .Z(n453) );
  GTECH_NOT U598 ( .A(n570), .Z(N105) );
  GTECH_AOI222 U599 ( .A(n374), .B(n457), .C(n376), .D(n458), .E(n456), .F(
        n372), .Z(n570) );
  GTECH_XOR2 U600 ( .A(n571), .B(n564), .Z(n456) );
  GTECH_ADD_ABC U601 ( .A(n40), .B(n360), .C(n572), .COUT(n564) );
  GTECH_NOT U602 ( .A(n573), .Z(n458) );
  GTECH_XOR2 U603 ( .A(n571), .B(n574), .Z(n573) );
  GTECH_NOT U604 ( .A(n569), .Z(n574) );
  GTECH_OAI21 U605 ( .A(n40), .B(n575), .C(n576), .Z(n569) );
  GTECH_OAI21 U606 ( .A(n360), .B(n461), .C(n577), .Z(n576) );
  GTECH_XOR2 U607 ( .A(n567), .B(n39), .Z(n571) );
  GTECH_NOT U608 ( .A(n361), .Z(n567) );
  GTECH_NOT U609 ( .A(n39), .Z(n457) );
  GTECH_NOT U610 ( .A(n578), .Z(N104) );
  GTECH_AOI222 U611 ( .A(n374), .B(n461), .C(n376), .D(n462), .E(n460), .F(
        n372), .Z(n578) );
  GTECH_XOR2 U612 ( .A(n579), .B(n572), .Z(n460) );
  GTECH_ADD_ABC U613 ( .A(n41), .B(n359), .C(n580), .COUT(n572) );
  GTECH_NOT U614 ( .A(n581), .Z(n462) );
  GTECH_XOR2 U615 ( .A(n579), .B(n582), .Z(n581) );
  GTECH_NOT U616 ( .A(n577), .Z(n582) );
  GTECH_OAI21 U617 ( .A(n41), .B(n583), .C(n584), .Z(n577) );
  GTECH_OAI21 U618 ( .A(n359), .B(n465), .C(n585), .Z(n584) );
  GTECH_XOR2 U619 ( .A(n575), .B(n40), .Z(n579) );
  GTECH_NOT U620 ( .A(n360), .Z(n575) );
  GTECH_NOT U621 ( .A(n40), .Z(n461) );
  GTECH_NOT U622 ( .A(n586), .Z(N103) );
  GTECH_AOI222 U623 ( .A(n374), .B(n465), .C(n376), .D(n466), .E(n464), .F(
        n372), .Z(n586) );
  GTECH_XOR2 U624 ( .A(n587), .B(n580), .Z(n464) );
  GTECH_ADD_ABC U625 ( .A(n42), .B(n358), .C(n588), .COUT(n580) );
  GTECH_NOT U626 ( .A(n589), .Z(n466) );
  GTECH_XOR2 U627 ( .A(n587), .B(n590), .Z(n589) );
  GTECH_NOT U628 ( .A(n585), .Z(n590) );
  GTECH_OAI21 U629 ( .A(n42), .B(n591), .C(n592), .Z(n585) );
  GTECH_OAI21 U630 ( .A(n358), .B(n470), .C(n593), .Z(n592) );
  GTECH_XOR2 U631 ( .A(n583), .B(n41), .Z(n587) );
  GTECH_NOT U632 ( .A(n359), .Z(n583) );
  GTECH_NOT U633 ( .A(n41), .Z(n465) );
  GTECH_NOT U634 ( .A(n594), .Z(N102) );
  GTECH_AOI222 U635 ( .A(n374), .B(n470), .C(n376), .D(n471), .E(n469), .F(
        n372), .Z(n594) );
  GTECH_XOR2 U636 ( .A(n595), .B(n588), .Z(n469) );
  GTECH_ADD_ABC U637 ( .A(n43), .B(n357), .C(n596), .COUT(n588) );
  GTECH_NOT U638 ( .A(n597), .Z(n471) );
  GTECH_XOR2 U639 ( .A(n595), .B(n598), .Z(n597) );
  GTECH_NOT U640 ( .A(n593), .Z(n598) );
  GTECH_OAI21 U641 ( .A(n43), .B(n599), .C(n600), .Z(n593) );
  GTECH_OAI21 U642 ( .A(n357), .B(n474), .C(n601), .Z(n600) );
  GTECH_XOR2 U643 ( .A(n591), .B(n42), .Z(n595) );
  GTECH_NOT U644 ( .A(n358), .Z(n591) );
  GTECH_NOT U645 ( .A(n42), .Z(n470) );
  GTECH_NOT U646 ( .A(n602), .Z(N101) );
  GTECH_AOI222 U647 ( .A(n374), .B(n474), .C(n376), .D(n475), .E(n473), .F(
        n372), .Z(n602) );
  GTECH_XOR2 U648 ( .A(n603), .B(n596), .Z(n473) );
  GTECH_ADD_ABC U649 ( .A(n356), .B(n29), .C(n604), .COUT(n596) );
  GTECH_NOT U650 ( .A(n605), .Z(n475) );
  GTECH_XOR2 U651 ( .A(n603), .B(n606), .Z(n605) );
  GTECH_NOT U652 ( .A(n601), .Z(n606) );
  GTECH_OAI21 U653 ( .A(n29), .B(n607), .C(n608), .Z(n601) );
  GTECH_OAI21 U654 ( .A(n356), .B(n478), .C(n609), .Z(n608) );
  GTECH_NOT U655 ( .A(n356), .Z(n607) );
  GTECH_XOR2 U656 ( .A(n599), .B(n43), .Z(n603) );
  GTECH_NOT U657 ( .A(n357), .Z(n599) );
  GTECH_NOT U658 ( .A(n43), .Z(n474) );
  GTECH_NOT U659 ( .A(n610), .Z(N100) );
  GTECH_AOI222 U660 ( .A(n477), .B(n372), .C(n374), .D(n478), .E(n376), .F(
        n479), .Z(n610) );
  GTECH_NOT U661 ( .A(n611), .Z(n479) );
  GTECH_XOR2 U662 ( .A(n612), .B(n613), .Z(n611) );
  GTECH_NOT U663 ( .A(n609), .Z(n613) );
  GTECH_OAI21 U664 ( .A(n11), .B(n614), .C(n615), .Z(n609) );
  GTECH_OAI21 U665 ( .A(n355), .B(n375), .C(n484), .Z(n615) );
  GTECH_NAND2 U666 ( .A(n12), .B(n490), .Z(n484) );
  GTECH_NOT U667 ( .A(n11), .Z(n375) );
  GTECH_NOT U668 ( .A(n355), .Z(n614) );
  GTECH_NOT U669 ( .A(n384), .Z(n376) );
  GTECH_NAND2 U670 ( .A(N82), .B(n10), .Z(n384) );
  GTECH_NOT U671 ( .A(n616), .Z(N82) );
  GTECH_NOT U672 ( .A(n617), .Z(n374) );
  GTECH_MUX2 U673 ( .A(n616), .B(n618), .S(n10), .Z(n617) );
  GTECH_NAND2 U674 ( .A(n28), .B(n385), .Z(n618) );
  GTECH_NAND2 U675 ( .A(n385), .B(n494), .Z(n616) );
  GTECH_NOT U676 ( .A(n28), .Z(n494) );
  GTECH_NOT U677 ( .A(n383), .Z(n372) );
  GTECH_NAND3 U678 ( .A(n385), .B(n492), .C(n28), .Z(n383) );
  GTECH_NOT U679 ( .A(n10), .Z(n492) );
  GTECH_NOT U680 ( .A(n407), .Z(n385) );
  GTECH_OAI21 U681 ( .A(n403), .B(n404), .C(n619), .Z(n407) );
  GTECH_AND2 U682 ( .A(n405), .B(n406), .Z(n619) );
  GTECH_NOT U683 ( .A(Rst), .Z(n406) );
  GTECH_NOT U684 ( .A(Ld), .Z(n405) );
  GTECH_NOT U685 ( .A(n9), .Z(n404) );
  GTECH_NAND2 U686 ( .A(n8), .B(n409), .Z(n403) );
  GTECH_NOT U687 ( .A(n412), .Z(n409) );
  GTECH_NAND2 U688 ( .A(n7), .B(n411), .Z(n412) );
  GTECH_NOT U689 ( .A(n620), .Z(n411) );
  GTECH_NAND2 U690 ( .A(n6), .B(n353), .Z(n620) );
  GTECH_XOR2 U691 ( .A(n612), .B(n604), .Z(n477) );
  GTECH_ADD_ABC U692 ( .A(n355), .B(n11), .C(n488), .COUT(n604) );
  GTECH_NAND2 U693 ( .A(n379), .B(n490), .Z(n488) );
  GTECH_NOT U694 ( .A(n354), .Z(n490) );
  GTECH_NOT U695 ( .A(n12), .Z(n379) );
  GTECH_XOR2 U696 ( .A(n478), .B(n356), .Z(n612) );
  GTECH_NOT U697 ( .A(n29), .Z(n478) );
endmodule

