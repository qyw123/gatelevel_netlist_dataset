
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366;

  GTECH_MUX2 U125 ( .A(n264), .B(n265), .S(n266), .Z(sum[9]) );
  GTECH_XOR2 U126 ( .A(n267), .B(n268), .Z(n265) );
  GTECH_XOR2 U127 ( .A(n269), .B(n268), .Z(n264) );
  GTECH_OA21 U128 ( .A(b[9]), .B(a[9]), .C(n270), .Z(n268) );
  GTECH_NOT U129 ( .A(n271), .Z(n270) );
  GTECH_XNOR2 U130 ( .A(n272), .B(n266), .Z(sum[8]) );
  GTECH_MUX2 U131 ( .A(n273), .B(n274), .S(n275), .Z(sum[7]) );
  GTECH_XNOR2 U132 ( .A(n276), .B(n277), .Z(n274) );
  GTECH_AOI21 U133 ( .A(n278), .B(n279), .C(n280), .Z(n277) );
  GTECH_XNOR2 U134 ( .A(n276), .B(n281), .Z(n273) );
  GTECH_XOR2 U135 ( .A(a[7]), .B(b[7]), .Z(n276) );
  GTECH_MUX2 U136 ( .A(n282), .B(n283), .S(n275), .Z(sum[6]) );
  GTECH_XOR2 U137 ( .A(n279), .B(n284), .Z(n283) );
  GTECH_OAI2N2 U138 ( .A(n285), .B(n286), .C(a[5]), .D(b[5]), .Z(n279) );
  GTECH_XOR2 U139 ( .A(n287), .B(n284), .Z(n282) );
  GTECH_AND_NOT U140 ( .A(n278), .B(n280), .Z(n284) );
  GTECH_MUX2 U141 ( .A(n288), .B(n289), .S(n275), .Z(sum[5]) );
  GTECH_XNOR2 U142 ( .A(n286), .B(n290), .Z(n289) );
  GTECH_XOR2 U143 ( .A(n291), .B(n290), .Z(n288) );
  GTECH_AOI21 U144 ( .A(b[5]), .B(a[5]), .C(n285), .Z(n290) );
  GTECH_NOT U145 ( .A(n292), .Z(n285) );
  GTECH_OR_NOT U146 ( .A(n293), .B(n294), .Z(sum[4]) );
  GTECH_AO21 U147 ( .A(n291), .B(n286), .C(n275), .Z(n294) );
  GTECH_MUX2 U148 ( .A(n295), .B(n296), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U149 ( .A(n297), .B(n298), .Z(n296) );
  GTECH_XOR2 U150 ( .A(n297), .B(n299), .Z(n295) );
  GTECH_AOI21 U151 ( .A(n300), .B(n301), .C(n302), .Z(n299) );
  GTECH_XNOR2 U152 ( .A(a[3]), .B(b[3]), .Z(n297) );
  GTECH_MUX2 U153 ( .A(n303), .B(n304), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U154 ( .A(n305), .B(n306), .Z(n304) );
  GTECH_XOR2 U155 ( .A(n301), .B(n306), .Z(n303) );
  GTECH_AND_NOT U156 ( .A(n300), .B(n302), .Z(n306) );
  GTECH_OR_NOT U157 ( .A(n307), .B(n308), .Z(n301) );
  GTECH_NAND3 U158 ( .A(b[0]), .B(n309), .C(a[0]), .Z(n308) );
  GTECH_MUX2 U159 ( .A(n310), .B(n311), .S(cin), .Z(sum[1]) );
  GTECH_XOR2 U160 ( .A(n312), .B(n313), .Z(n311) );
  GTECH_XOR2 U161 ( .A(n312), .B(n314), .Z(n310) );
  GTECH_AND2 U162 ( .A(a[0]), .B(b[0]), .Z(n314) );
  GTECH_AND_NOT U163 ( .A(n309), .B(n307), .Z(n312) );
  GTECH_MUX2 U164 ( .A(n315), .B(n316), .S(n317), .Z(sum[15]) );
  GTECH_XOR2 U165 ( .A(n318), .B(n319), .Z(n316) );
  GTECH_XOR2 U166 ( .A(n318), .B(n320), .Z(n315) );
  GTECH_OA21 U167 ( .A(n321), .B(n322), .C(n323), .Z(n320) );
  GTECH_XNOR2 U168 ( .A(n324), .B(n325), .Z(n318) );
  GTECH_MUX2 U169 ( .A(n326), .B(n327), .S(n317), .Z(sum[14]) );
  GTECH_XOR2 U170 ( .A(n328), .B(n329), .Z(n327) );
  GTECH_XOR2 U171 ( .A(n328), .B(n322), .Z(n326) );
  GTECH_AOI21 U172 ( .A(n330), .B(n331), .C(n332), .Z(n322) );
  GTECH_OR_NOT U173 ( .A(n321), .B(n323), .Z(n328) );
  GTECH_MUX2 U174 ( .A(n333), .B(n334), .S(n335), .Z(sum[13]) );
  GTECH_OA21 U175 ( .A(n330), .B(n317), .C(n336), .Z(n335) );
  GTECH_OR_NOT U176 ( .A(n332), .B(n331), .Z(n334) );
  GTECH_XOR2 U177 ( .A(b[13]), .B(a[13]), .Z(n333) );
  GTECH_OR_NOT U178 ( .A(n337), .B(n338), .Z(sum[12]) );
  GTECH_AO21 U179 ( .A(n336), .B(n339), .C(n340), .Z(n338) );
  GTECH_MUX2 U180 ( .A(n341), .B(n342), .S(n266), .Z(sum[11]) );
  GTECH_XOR2 U181 ( .A(n343), .B(n344), .Z(n342) );
  GTECH_AOI21 U182 ( .A(n345), .B(n346), .C(n347), .Z(n344) );
  GTECH_XNOR2 U183 ( .A(n343), .B(n348), .Z(n341) );
  GTECH_XNOR2 U184 ( .A(a[11]), .B(b[11]), .Z(n343) );
  GTECH_MUX2 U185 ( .A(n349), .B(n350), .S(n266), .Z(sum[10]) );
  GTECH_XNOR2 U186 ( .A(n351), .B(n346), .Z(n350) );
  GTECH_OA21 U187 ( .A(n267), .B(n271), .C(n352), .Z(n346) );
  GTECH_XNOR2 U188 ( .A(n351), .B(n353), .Z(n349) );
  GTECH_OR_NOT U189 ( .A(n347), .B(n345), .Z(n351) );
  GTECH_XNOR2 U190 ( .A(cin), .B(n354), .Z(sum[0]) );
  GTECH_AO21 U191 ( .A(n317), .B(n355), .C(n337), .Z(cout) );
  GTECH_AND3 U192 ( .A(n336), .B(n339), .C(n340), .Z(n337) );
  GTECH_NOT U193 ( .A(n317), .Z(n340) );
  GTECH_NOT U194 ( .A(n330), .Z(n339) );
  GTECH_AND2 U195 ( .A(b[12]), .B(a[12]), .Z(n330) );
  GTECH_OAI22 U196 ( .A(n319), .B(n324), .C(n356), .D(n325), .Z(n355) );
  GTECH_NOT U197 ( .A(b[15]), .Z(n325) );
  GTECH_AND_NOT U198 ( .A(n319), .B(a[15]), .Z(n356) );
  GTECH_NOT U199 ( .A(a[15]), .Z(n324) );
  GTECH_OA21 U200 ( .A(n321), .B(n329), .C(n323), .Z(n319) );
  GTECH_NAND2 U201 ( .A(b[14]), .B(a[14]), .Z(n323) );
  GTECH_AOI21 U202 ( .A(n336), .B(n331), .C(n332), .Z(n329) );
  GTECH_AND_NOT U203 ( .A(b[13]), .B(n357), .Z(n332) );
  GTECH_NOT U204 ( .A(a[13]), .Z(n357) );
  GTECH_OR2 U205 ( .A(b[13]), .B(a[13]), .Z(n331) );
  GTECH_OR2 U206 ( .A(b[12]), .B(a[12]), .Z(n336) );
  GTECH_NOT U207 ( .A(n358), .Z(n321) );
  GTECH_OR2 U208 ( .A(a[14]), .B(b[14]), .Z(n358) );
  GTECH_MUX2 U209 ( .A(n359), .B(n272), .S(n266), .Z(n317) );
  GTECH_AOI21 U210 ( .A(n360), .B(n361), .C(n293), .Z(n266) );
  GTECH_AND3 U211 ( .A(n291), .B(n286), .C(n275), .Z(n293) );
  GTECH_NAND2 U212 ( .A(b[4]), .B(a[4]), .Z(n286) );
  GTECH_OAI2N2 U213 ( .A(n281), .B(n362), .C(n363), .D(b[7]), .Z(n361) );
  GTECH_OR_NOT U214 ( .A(a[7]), .B(n281), .Z(n363) );
  GTECH_NOT U215 ( .A(a[7]), .Z(n362) );
  GTECH_AOI21 U216 ( .A(n278), .B(n287), .C(n280), .Z(n281) );
  GTECH_AND2 U217 ( .A(b[6]), .B(a[6]), .Z(n280) );
  GTECH_AO22 U218 ( .A(n291), .B(n292), .C(a[5]), .D(b[5]), .Z(n287) );
  GTECH_OR2 U219 ( .A(a[5]), .B(b[5]), .Z(n292) );
  GTECH_OR2 U220 ( .A(a[4]), .B(b[4]), .Z(n291) );
  GTECH_OR2 U221 ( .A(b[6]), .B(a[6]), .Z(n278) );
  GTECH_NOT U222 ( .A(n275), .Z(n360) );
  GTECH_MUX2 U223 ( .A(n354), .B(n364), .S(cin), .Z(n275) );
  GTECH_AOI21 U224 ( .A(n298), .B(a[3]), .C(n365), .Z(n364) );
  GTECH_OA21 U225 ( .A(n298), .B(a[3]), .C(b[3]), .Z(n365) );
  GTECH_AO21 U226 ( .A(n300), .B(n305), .C(n302), .Z(n298) );
  GTECH_AND2 U227 ( .A(b[2]), .B(a[2]), .Z(n302) );
  GTECH_AO21 U228 ( .A(n309), .B(n313), .C(n307), .Z(n305) );
  GTECH_AND2 U229 ( .A(b[1]), .B(a[1]), .Z(n307) );
  GTECH_OR2 U230 ( .A(a[0]), .B(b[0]), .Z(n313) );
  GTECH_OR2 U231 ( .A(a[1]), .B(b[1]), .Z(n309) );
  GTECH_OR2 U232 ( .A(b[2]), .B(a[2]), .Z(n300) );
  GTECH_XNOR2 U233 ( .A(a[0]), .B(b[0]), .Z(n354) );
  GTECH_AND_NOT U234 ( .A(n269), .B(n267), .Z(n272) );
  GTECH_AND2 U235 ( .A(a[8]), .B(b[8]), .Z(n267) );
  GTECH_OA21 U236 ( .A(a[11]), .B(n348), .C(n366), .Z(n359) );
  GTECH_AO21 U237 ( .A(a[11]), .B(n348), .C(b[11]), .Z(n366) );
  GTECH_AO21 U238 ( .A(n353), .B(n345), .C(n347), .Z(n348) );
  GTECH_AND2 U239 ( .A(b[10]), .B(a[10]), .Z(n347) );
  GTECH_OR2 U240 ( .A(a[10]), .B(b[10]), .Z(n345) );
  GTECH_OA21 U241 ( .A(n269), .B(n271), .C(n352), .Z(n353) );
  GTECH_OR2 U242 ( .A(a[9]), .B(b[9]), .Z(n352) );
  GTECH_AND2 U243 ( .A(b[9]), .B(a[9]), .Z(n271) );
  GTECH_OR2 U244 ( .A(a[8]), .B(b[8]), .Z(n269) );
endmodule

