
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375;

  GTECH_OAI22 U133 ( .A(n272), .B(n273), .C(n274), .D(n275), .Z(sum[9]) );
  GTECH_XOR2 U134 ( .A(n276), .B(n277), .Z(n274) );
  GTECH_XNOR2 U135 ( .A(n278), .B(n277), .Z(n273) );
  GTECH_AND_NOT U136 ( .A(n279), .B(n280), .Z(n277) );
  GTECH_NAND2 U137 ( .A(n281), .B(n282), .Z(sum[8]) );
  GTECH_OAI21 U138 ( .A(n278), .B(n276), .C(n272), .Z(n281) );
  GTECH_OAI22 U139 ( .A(n283), .B(n284), .C(n285), .D(n286), .Z(sum[7]) );
  GTECH_XNOR2 U140 ( .A(n287), .B(n288), .Z(n285) );
  GTECH_XNOR2 U141 ( .A(n288), .B(n289), .Z(n284) );
  GTECH_OA21 U142 ( .A(a[6]), .B(n290), .C(n291), .Z(n289) );
  GTECH_AO21 U143 ( .A(n290), .B(a[6]), .C(b[6]), .Z(n291) );
  GTECH_XOR2 U144 ( .A(a[7]), .B(b[7]), .Z(n288) );
  GTECH_OAI22 U145 ( .A(n292), .B(n283), .C(n293), .D(n286), .Z(sum[6]) );
  GTECH_XNOR2 U146 ( .A(n294), .B(n295), .Z(n293) );
  GTECH_XNOR2 U147 ( .A(n290), .B(n295), .Z(n292) );
  GTECH_XOR2 U148 ( .A(a[6]), .B(b[6]), .Z(n295) );
  GTECH_AO21 U149 ( .A(n296), .B(n297), .C(n298), .Z(n290) );
  GTECH_OAI2N2 U150 ( .A(n299), .B(n300), .C(n301), .D(n299), .Z(sum[5]) );
  GTECH_OAI21 U151 ( .A(n297), .B(n283), .C(n302), .Z(n301) );
  GTECH_AOI21 U152 ( .A(n302), .B(n283), .C(n297), .Z(n300) );
  GTECH_NOT U153 ( .A(n286), .Z(n283) );
  GTECH_NOR2 U154 ( .A(n303), .B(n298), .Z(n299) );
  GTECH_XNOR2 U155 ( .A(n286), .B(n304), .Z(sum[4]) );
  GTECH_OAI22 U156 ( .A(n305), .B(n306), .C(cin), .D(n307), .Z(sum[3]) );
  GTECH_XOR2 U157 ( .A(n308), .B(n309), .Z(n307) );
  GTECH_OA21 U158 ( .A(n310), .B(n311), .C(n312), .Z(n308) );
  GTECH_XNOR2 U159 ( .A(n313), .B(n309), .Z(n306) );
  GTECH_XOR2 U160 ( .A(a[3]), .B(b[3]), .Z(n309) );
  GTECH_OAI22 U161 ( .A(n305), .B(n314), .C(cin), .D(n315), .Z(sum[2]) );
  GTECH_XOR2 U162 ( .A(n316), .B(n311), .Z(n315) );
  GTECH_AOI21 U163 ( .A(n317), .B(n318), .C(n319), .Z(n311) );
  GTECH_XOR2 U164 ( .A(n316), .B(n320), .Z(n314) );
  GTECH_AND_NOT U165 ( .A(n312), .B(n310), .Z(n316) );
  GTECH_OAI2N2 U166 ( .A(n321), .B(n322), .C(n323), .D(n321), .Z(sum[1]) );
  GTECH_OAI21 U167 ( .A(cin), .B(n318), .C(n324), .Z(n323) );
  GTECH_AOI21 U168 ( .A(n324), .B(cin), .C(n318), .Z(n322) );
  GTECH_AND2 U169 ( .A(b[0]), .B(a[0]), .Z(n318) );
  GTECH_NOR2 U170 ( .A(n325), .B(n319), .Z(n321) );
  GTECH_OAI22 U171 ( .A(n326), .B(n327), .C(n328), .D(n329), .Z(sum[15]) );
  GTECH_XNOR2 U172 ( .A(n330), .B(n331), .Z(n329) );
  GTECH_XOR2 U173 ( .A(n332), .B(n331), .Z(n327) );
  GTECH_XOR2 U174 ( .A(a[15]), .B(b[15]), .Z(n331) );
  GTECH_AOI21 U175 ( .A(n333), .B(n334), .C(n335), .Z(n332) );
  GTECH_OAI22 U176 ( .A(n326), .B(n336), .C(n328), .D(n337), .Z(sum[14]) );
  GTECH_XNOR2 U177 ( .A(n338), .B(n339), .Z(n337) );
  GTECH_XNOR2 U178 ( .A(n334), .B(n339), .Z(n336) );
  GTECH_AND_NOT U179 ( .A(n333), .B(n335), .Z(n339) );
  GTECH_AOI21 U180 ( .A(n340), .B(n341), .C(n342), .Z(n334) );
  GTECH_OAI22 U181 ( .A(n326), .B(n343), .C(n328), .D(n344), .Z(sum[13]) );
  GTECH_XOR2 U182 ( .A(n345), .B(n346), .Z(n344) );
  GTECH_XNOR2 U183 ( .A(n341), .B(n346), .Z(n343) );
  GTECH_OAI21 U184 ( .A(a[13]), .B(b[13]), .C(n340), .Z(n346) );
  GTECH_NAND2 U185 ( .A(n347), .B(n348), .Z(sum[12]) );
  GTECH_AO21 U186 ( .A(n341), .B(n345), .C(n328), .Z(n347) );
  GTECH_OAI22 U187 ( .A(n349), .B(n272), .C(n350), .D(n275), .Z(sum[11]) );
  GTECH_XNOR2 U188 ( .A(n351), .B(n352), .Z(n350) );
  GTECH_XOR2 U189 ( .A(n353), .B(n352), .Z(n349) );
  GTECH_XOR2 U190 ( .A(a[11]), .B(b[11]), .Z(n352) );
  GTECH_OA21 U191 ( .A(n354), .B(n355), .C(n356), .Z(n353) );
  GTECH_OAI22 U192 ( .A(n357), .B(n272), .C(n358), .D(n275), .Z(sum[10]) );
  GTECH_XOR2 U193 ( .A(n359), .B(n360), .Z(n358) );
  GTECH_XOR2 U194 ( .A(n359), .B(n355), .Z(n357) );
  GTECH_OA21 U195 ( .A(n280), .B(n361), .C(n279), .Z(n355) );
  GTECH_NOT U196 ( .A(n278), .Z(n361) );
  GTECH_AND_NOT U197 ( .A(n356), .B(n354), .Z(n359) );
  GTECH_XNOR2 U198 ( .A(n305), .B(n362), .Z(sum[0]) );
  GTECH_OAI21 U199 ( .A(n328), .B(n363), .C(n348), .Z(cout) );
  GTECH_NAND3 U200 ( .A(n341), .B(n345), .C(n328), .Z(n348) );
  GTECH_NOT U201 ( .A(n364), .Z(n345) );
  GTECH_NAND2 U202 ( .A(b[12]), .B(a[12]), .Z(n341) );
  GTECH_AOI21 U203 ( .A(n330), .B(a[15]), .C(n365), .Z(n363) );
  GTECH_OA21 U204 ( .A(a[15]), .B(n330), .C(b[15]), .Z(n365) );
  GTECH_AO21 U205 ( .A(n333), .B(n338), .C(n335), .Z(n330) );
  GTECH_AND2 U206 ( .A(a[14]), .B(b[14]), .Z(n335) );
  GTECH_AOI21 U207 ( .A(n340), .B(n364), .C(n342), .Z(n338) );
  GTECH_NOR2 U208 ( .A(b[13]), .B(a[13]), .Z(n342) );
  GTECH_NOR2 U209 ( .A(b[12]), .B(a[12]), .Z(n364) );
  GTECH_NAND2 U210 ( .A(a[13]), .B(b[13]), .Z(n340) );
  GTECH_NOT U211 ( .A(n366), .Z(n333) );
  GTECH_NOR2 U212 ( .A(a[14]), .B(b[14]), .Z(n366) );
  GTECH_NOT U213 ( .A(n326), .Z(n328) );
  GTECH_OAI21 U214 ( .A(n367), .B(n275), .C(n282), .Z(n326) );
  GTECH_OR3 U215 ( .A(n278), .B(n276), .C(n272), .Z(n282) );
  GTECH_NOT U216 ( .A(n275), .Z(n272) );
  GTECH_AND2 U217 ( .A(b[8]), .B(a[8]), .Z(n278) );
  GTECH_AOI2N2 U218 ( .A(n286), .B(n304), .C(n368), .D(n286), .Z(n275) );
  GTECH_AOI21 U219 ( .A(n287), .B(a[7]), .C(n369), .Z(n368) );
  GTECH_OA21 U220 ( .A(a[7]), .B(n287), .C(b[7]), .Z(n369) );
  GTECH_AO21 U221 ( .A(n294), .B(a[6]), .C(n370), .Z(n287) );
  GTECH_OA21 U222 ( .A(a[6]), .B(n294), .C(b[6]), .Z(n370) );
  GTECH_AO21 U223 ( .A(n302), .B(n296), .C(n298), .Z(n294) );
  GTECH_AND2 U224 ( .A(a[5]), .B(b[5]), .Z(n298) );
  GTECH_NOT U225 ( .A(n303), .Z(n296) );
  GTECH_NOR2 U226 ( .A(a[5]), .B(b[5]), .Z(n303) );
  GTECH_AND_NOT U227 ( .A(n302), .B(n297), .Z(n304) );
  GTECH_AND2 U228 ( .A(a[4]), .B(b[4]), .Z(n297) );
  GTECH_NOT U229 ( .A(n371), .Z(n302) );
  GTECH_NOR2 U230 ( .A(a[4]), .B(b[4]), .Z(n371) );
  GTECH_AOI2N2 U231 ( .A(n305), .B(n362), .C(n372), .D(n305), .Z(n286) );
  GTECH_AOI21 U232 ( .A(n313), .B(a[3]), .C(n373), .Z(n372) );
  GTECH_OA21 U233 ( .A(a[3]), .B(n313), .C(b[3]), .Z(n373) );
  GTECH_OAI21 U234 ( .A(n320), .B(n310), .C(n312), .Z(n313) );
  GTECH_NAND2 U235 ( .A(a[2]), .B(b[2]), .Z(n312) );
  GTECH_NOR2 U236 ( .A(a[2]), .B(b[2]), .Z(n310) );
  GTECH_AOI21 U237 ( .A(n317), .B(n324), .C(n319), .Z(n320) );
  GTECH_AND2 U238 ( .A(a[1]), .B(b[1]), .Z(n319) );
  GTECH_NOT U239 ( .A(n374), .Z(n324) );
  GTECH_NOR2 U240 ( .A(b[0]), .B(a[0]), .Z(n374) );
  GTECH_NOT U241 ( .A(n325), .Z(n317) );
  GTECH_NOR2 U242 ( .A(a[1]), .B(b[1]), .Z(n325) );
  GTECH_XOR2 U243 ( .A(a[0]), .B(b[0]), .Z(n362) );
  GTECH_NOT U244 ( .A(cin), .Z(n305) );
  GTECH_AOI21 U245 ( .A(n351), .B(a[11]), .C(n375), .Z(n367) );
  GTECH_OA21 U246 ( .A(a[11]), .B(n351), .C(b[11]), .Z(n375) );
  GTECH_OAI21 U247 ( .A(n360), .B(n354), .C(n356), .Z(n351) );
  GTECH_NAND2 U248 ( .A(a[10]), .B(b[10]), .Z(n356) );
  GTECH_NOR2 U249 ( .A(a[10]), .B(b[10]), .Z(n354) );
  GTECH_OA21 U250 ( .A(n276), .B(n280), .C(n279), .Z(n360) );
  GTECH_NAND2 U251 ( .A(a[9]), .B(b[9]), .Z(n279) );
  GTECH_NOR2 U252 ( .A(a[9]), .B(b[9]), .Z(n280) );
  GTECH_NOR2 U253 ( .A(b[8]), .B(a[8]), .Z(n276) );
endmodule

