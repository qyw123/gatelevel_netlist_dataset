
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378;

  GTECH_MUX2 U136 ( .A(n275), .B(n276), .S(n277), .Z(sum[9]) );
  GTECH_XNOR2 U137 ( .A(n278), .B(n279), .Z(n276) );
  GTECH_XNOR2 U138 ( .A(n280), .B(n278), .Z(n275) );
  GTECH_OAI21 U139 ( .A(a[9]), .B(b[9]), .C(n281), .Z(n278) );
  GTECH_NOT U140 ( .A(n282), .Z(n281) );
  GTECH_OAI21 U141 ( .A(n283), .B(n284), .C(n285), .Z(sum[8]) );
  GTECH_NOR2 U142 ( .A(n286), .B(n280), .Z(n283) );
  GTECH_MUX2 U143 ( .A(n287), .B(n288), .S(n289), .Z(sum[7]) );
  GTECH_XNOR2 U144 ( .A(n290), .B(n291), .Z(n288) );
  GTECH_XOR2 U145 ( .A(n290), .B(n292), .Z(n287) );
  GTECH_OA21 U146 ( .A(n293), .B(n294), .C(n295), .Z(n292) );
  GTECH_XNOR2 U147 ( .A(a[7]), .B(b[7]), .Z(n290) );
  GTECH_MUX2 U148 ( .A(n296), .B(n297), .S(n289), .Z(sum[6]) );
  GTECH_XOR2 U149 ( .A(n298), .B(n299), .Z(n297) );
  GTECH_XOR2 U150 ( .A(n298), .B(n294), .Z(n296) );
  GTECH_OA21 U151 ( .A(n300), .B(n301), .C(n302), .Z(n294) );
  GTECH_OR2 U152 ( .A(n293), .B(n303), .Z(n298) );
  GTECH_MUX2 U153 ( .A(n304), .B(n305), .S(n306), .Z(sum[5]) );
  GTECH_NOR2 U154 ( .A(n307), .B(n300), .Z(n306) );
  GTECH_OAI2N2 U155 ( .A(b[4]), .B(a[4]), .C(n301), .D(n308), .Z(n305) );
  GTECH_OR_NOT U156 ( .A(n309), .B(b[4]), .Z(n301) );
  GTECH_OAI21 U157 ( .A(n308), .B(n309), .C(n310), .Z(n304) );
  GTECH_OAI21 U158 ( .A(a[4]), .B(n289), .C(b[4]), .Z(n310) );
  GTECH_XNOR2 U159 ( .A(n311), .B(n308), .Z(sum[4]) );
  GTECH_NOT U160 ( .A(n289), .Z(n308) );
  GTECH_MUX2 U161 ( .A(n312), .B(n313), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U162 ( .A(n314), .B(n315), .Z(n313) );
  GTECH_XOR2 U163 ( .A(n314), .B(n316), .Z(n312) );
  GTECH_OA21 U164 ( .A(n317), .B(n318), .C(n319), .Z(n316) );
  GTECH_XNOR2 U165 ( .A(a[3]), .B(b[3]), .Z(n314) );
  GTECH_MUX2 U166 ( .A(n320), .B(n321), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U167 ( .A(n322), .B(n323), .Z(n321) );
  GTECH_XNOR2 U168 ( .A(n318), .B(n322), .Z(n320) );
  GTECH_NOR2 U169 ( .A(n324), .B(n317), .Z(n322) );
  GTECH_AOI21 U170 ( .A(n325), .B(n326), .C(n327), .Z(n318) );
  GTECH_MUX2 U171 ( .A(n328), .B(n329), .S(n330), .Z(sum[1]) );
  GTECH_AND_NOT U172 ( .A(n325), .B(n327), .Z(n330) );
  GTECH_OAI21 U173 ( .A(cin), .B(n326), .C(n331), .Z(n329) );
  GTECH_AO21 U174 ( .A(n331), .B(cin), .C(n326), .Z(n328) );
  GTECH_AND2 U175 ( .A(a[0]), .B(b[0]), .Z(n326) );
  GTECH_MUX2 U176 ( .A(n332), .B(n333), .S(n334), .Z(sum[15]) );
  GTECH_XOR2 U177 ( .A(n335), .B(n336), .Z(n333) );
  GTECH_AOI21 U178 ( .A(n337), .B(n338), .C(n339), .Z(n336) );
  GTECH_XNOR2 U179 ( .A(n335), .B(n340), .Z(n332) );
  GTECH_XNOR2 U180 ( .A(a[15]), .B(b[15]), .Z(n335) );
  GTECH_MUX2 U181 ( .A(n341), .B(n342), .S(n334), .Z(sum[14]) );
  GTECH_XNOR2 U182 ( .A(n343), .B(n338), .Z(n342) );
  GTECH_OA21 U183 ( .A(n344), .B(n345), .C(n346), .Z(n338) );
  GTECH_XNOR2 U184 ( .A(n343), .B(n347), .Z(n341) );
  GTECH_OR_NOT U185 ( .A(n339), .B(n337), .Z(n343) );
  GTECH_MUX2 U186 ( .A(n348), .B(n349), .S(n334), .Z(sum[13]) );
  GTECH_XNOR2 U187 ( .A(n345), .B(n350), .Z(n349) );
  GTECH_XNOR2 U188 ( .A(n350), .B(n351), .Z(n348) );
  GTECH_OAI21 U189 ( .A(a[13]), .B(b[13]), .C(n352), .Z(n350) );
  GTECH_NOT U190 ( .A(n344), .Z(n352) );
  GTECH_OAI21 U191 ( .A(n334), .B(n353), .C(n354), .Z(sum[12]) );
  GTECH_AND_NOT U192 ( .A(n351), .B(n345), .Z(n353) );
  GTECH_MUX2 U193 ( .A(n355), .B(n356), .S(n277), .Z(sum[11]) );
  GTECH_XNOR2 U194 ( .A(n357), .B(n358), .Z(n356) );
  GTECH_XOR2 U195 ( .A(n357), .B(n359), .Z(n355) );
  GTECH_AOI21 U196 ( .A(n360), .B(n361), .C(n362), .Z(n359) );
  GTECH_XNOR2 U197 ( .A(a[11]), .B(b[11]), .Z(n357) );
  GTECH_MUX2 U198 ( .A(n363), .B(n364), .S(n277), .Z(sum[10]) );
  GTECH_XOR2 U199 ( .A(n365), .B(n366), .Z(n364) );
  GTECH_XOR2 U200 ( .A(n365), .B(n361), .Z(n363) );
  GTECH_OA21 U201 ( .A(n282), .B(n280), .C(n367), .Z(n361) );
  GTECH_AND_NOT U202 ( .A(n360), .B(n362), .Z(n365) );
  GTECH_XOR2 U203 ( .A(cin), .B(n368), .Z(sum[0]) );
  GTECH_OAI21 U204 ( .A(n334), .B(n369), .C(n354), .Z(cout) );
  GTECH_NAND3 U205 ( .A(n370), .B(n351), .C(n334), .Z(n354) );
  GTECH_NOT U206 ( .A(n345), .Z(n370) );
  GTECH_AND2 U207 ( .A(b[12]), .B(a[12]), .Z(n345) );
  GTECH_AOI21 U208 ( .A(n340), .B(a[15]), .C(n371), .Z(n369) );
  GTECH_OA21 U209 ( .A(a[15]), .B(n340), .C(b[15]), .Z(n371) );
  GTECH_AO21 U210 ( .A(n337), .B(n347), .C(n339), .Z(n340) );
  GTECH_AND2 U211 ( .A(b[14]), .B(a[14]), .Z(n339) );
  GTECH_OA21 U212 ( .A(n344), .B(n351), .C(n346), .Z(n347) );
  GTECH_OR2 U213 ( .A(a[13]), .B(b[13]), .Z(n346) );
  GTECH_OR2 U214 ( .A(a[12]), .B(b[12]), .Z(n351) );
  GTECH_AND2 U215 ( .A(b[13]), .B(a[13]), .Z(n344) );
  GTECH_OR2 U216 ( .A(a[14]), .B(b[14]), .Z(n337) );
  GTECH_OA21 U217 ( .A(n372), .B(n284), .C(n285), .Z(n334) );
  GTECH_OR3 U218 ( .A(n280), .B(n286), .C(n277), .Z(n285) );
  GTECH_NOT U219 ( .A(n279), .Z(n286) );
  GTECH_AND2 U220 ( .A(b[8]), .B(a[8]), .Z(n280) );
  GTECH_NOT U221 ( .A(n277), .Z(n284) );
  GTECH_MUX2 U222 ( .A(n311), .B(n373), .S(n289), .Z(n277) );
  GTECH_MUX2 U223 ( .A(n368), .B(n374), .S(cin), .Z(n289) );
  GTECH_OA21 U224 ( .A(a[3]), .B(n315), .C(n375), .Z(n374) );
  GTECH_AO21 U225 ( .A(n315), .B(a[3]), .C(b[3]), .Z(n375) );
  GTECH_OAI21 U226 ( .A(n323), .B(n317), .C(n319), .Z(n315) );
  GTECH_NOT U227 ( .A(n324), .Z(n319) );
  GTECH_AND2 U228 ( .A(b[2]), .B(a[2]), .Z(n324) );
  GTECH_NOR2 U229 ( .A(b[2]), .B(a[2]), .Z(n317) );
  GTECH_AOI21 U230 ( .A(n331), .B(n325), .C(n327), .Z(n323) );
  GTECH_AND2 U231 ( .A(a[1]), .B(b[1]), .Z(n327) );
  GTECH_OR2 U232 ( .A(a[1]), .B(b[1]), .Z(n325) );
  GTECH_OR2 U233 ( .A(b[0]), .B(a[0]), .Z(n331) );
  GTECH_XOR2 U234 ( .A(a[0]), .B(b[0]), .Z(n368) );
  GTECH_OA21 U235 ( .A(a[7]), .B(n291), .C(n376), .Z(n373) );
  GTECH_AO21 U236 ( .A(n291), .B(a[7]), .C(b[7]), .Z(n376) );
  GTECH_OAI21 U237 ( .A(n299), .B(n293), .C(n295), .Z(n291) );
  GTECH_NOT U238 ( .A(n303), .Z(n295) );
  GTECH_AND2 U239 ( .A(b[6]), .B(a[6]), .Z(n303) );
  GTECH_NOR2 U240 ( .A(b[6]), .B(a[6]), .Z(n293) );
  GTECH_OA21 U241 ( .A(n377), .B(n300), .C(n302), .Z(n299) );
  GTECH_NOT U242 ( .A(n307), .Z(n302) );
  GTECH_AND2 U243 ( .A(a[5]), .B(b[5]), .Z(n307) );
  GTECH_NOR2 U244 ( .A(a[5]), .B(b[5]), .Z(n300) );
  GTECH_AND_NOT U245 ( .A(n309), .B(b[4]), .Z(n377) );
  GTECH_NOT U246 ( .A(a[4]), .Z(n309) );
  GTECH_XOR2 U247 ( .A(a[4]), .B(b[4]), .Z(n311) );
  GTECH_AOI21 U248 ( .A(n358), .B(a[11]), .C(n378), .Z(n372) );
  GTECH_OA21 U249 ( .A(a[11]), .B(n358), .C(b[11]), .Z(n378) );
  GTECH_AO21 U250 ( .A(n360), .B(n366), .C(n362), .Z(n358) );
  GTECH_AND2 U251 ( .A(b[10]), .B(a[10]), .Z(n362) );
  GTECH_OA21 U252 ( .A(n282), .B(n279), .C(n367), .Z(n366) );
  GTECH_OR2 U253 ( .A(a[9]), .B(b[9]), .Z(n367) );
  GTECH_OR2 U254 ( .A(a[8]), .B(b[8]), .Z(n279) );
  GTECH_AND2 U255 ( .A(a[9]), .B(b[9]), .Z(n282) );
  GTECH_OR2 U256 ( .A(a[10]), .B(b[10]), .Z(n360) );
endmodule

