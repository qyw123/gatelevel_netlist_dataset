
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388;

  GTECH_MUX2 U138 ( .A(n277), .B(n278), .S(n279), .Z(sum[9]) );
  GTECH_XNOR2 U139 ( .A(n280), .B(n281), .Z(n278) );
  GTECH_XNOR2 U140 ( .A(n280), .B(n282), .Z(n277) );
  GTECH_AOI21 U141 ( .A(a[9]), .B(b[9]), .C(n283), .Z(n280) );
  GTECH_XNOR2 U142 ( .A(n279), .B(n284), .Z(sum[8]) );
  GTECH_MUX2 U143 ( .A(n285), .B(n286), .S(n287), .Z(sum[7]) );
  GTECH_XNOR2 U144 ( .A(n288), .B(n289), .Z(n286) );
  GTECH_AND_NOT U145 ( .A(n290), .B(n291), .Z(n289) );
  GTECH_OAI21 U146 ( .A(b[6]), .B(a[6]), .C(n292), .Z(n290) );
  GTECH_XOR2 U147 ( .A(n288), .B(n293), .Z(n285) );
  GTECH_XOR2 U148 ( .A(a[7]), .B(b[7]), .Z(n288) );
  GTECH_AO21 U149 ( .A(n294), .B(n291), .C(n295), .Z(sum[6]) );
  GTECH_NOT U150 ( .A(n296), .Z(n295) );
  GTECH_MUX2 U151 ( .A(n297), .B(n298), .S(b[6]), .Z(n296) );
  GTECH_OR2 U152 ( .A(n294), .B(a[6]), .Z(n298) );
  GTECH_XOR2 U153 ( .A(n299), .B(n294), .Z(n297) );
  GTECH_AO21 U154 ( .A(n300), .B(n301), .C(n292), .Z(n294) );
  GTECH_OAI21 U155 ( .A(n302), .B(n303), .C(n304), .Z(n292) );
  GTECH_OR2 U156 ( .A(n305), .B(n306), .Z(n303) );
  GTECH_MUX2 U157 ( .A(n307), .B(n308), .S(n309), .Z(sum[5]) );
  GTECH_AND_NOT U158 ( .A(n304), .B(n305), .Z(n309) );
  GTECH_OAI21 U159 ( .A(a[4]), .B(n301), .C(n310), .Z(n308) );
  GTECH_AO21 U160 ( .A(n301), .B(a[4]), .C(b[4]), .Z(n310) );
  GTECH_OAI2N2 U161 ( .A(n311), .B(n287), .C(b[4]), .D(a[4]), .Z(n307) );
  GTECH_XNOR2 U162 ( .A(n312), .B(n287), .Z(sum[4]) );
  GTECH_MUX2 U163 ( .A(n313), .B(n314), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U164 ( .A(n315), .B(n316), .Z(n314) );
  GTECH_XOR2 U165 ( .A(n317), .B(n315), .Z(n313) );
  GTECH_XOR2 U166 ( .A(a[3]), .B(b[3]), .Z(n315) );
  GTECH_OA21 U167 ( .A(a[2]), .B(n318), .C(n319), .Z(n317) );
  GTECH_AO21 U168 ( .A(n318), .B(a[2]), .C(b[2]), .Z(n319) );
  GTECH_MUX2 U169 ( .A(n320), .B(n321), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U170 ( .A(n322), .B(n323), .Z(n321) );
  GTECH_XNOR2 U171 ( .A(n322), .B(n318), .Z(n320) );
  GTECH_AO21 U172 ( .A(n324), .B(n325), .C(n326), .Z(n318) );
  GTECH_XNOR2 U173 ( .A(a[2]), .B(b[2]), .Z(n322) );
  GTECH_MUX2 U174 ( .A(n327), .B(n328), .S(n329), .Z(sum[1]) );
  GTECH_AND_NOT U175 ( .A(n324), .B(n326), .Z(n329) );
  GTECH_AO21 U176 ( .A(n330), .B(n331), .C(n332), .Z(n328) );
  GTECH_NOT U177 ( .A(cin), .Z(n330) );
  GTECH_AO21 U178 ( .A(n333), .B(cin), .C(n325), .Z(n327) );
  GTECH_MUX2 U179 ( .A(n334), .B(n335), .S(n336), .Z(sum[15]) );
  GTECH_XNOR2 U180 ( .A(n337), .B(n338), .Z(n335) );
  GTECH_XOR2 U181 ( .A(n337), .B(n339), .Z(n334) );
  GTECH_AND_NOT U182 ( .A(n340), .B(n341), .Z(n339) );
  GTECH_OAI21 U183 ( .A(b[14]), .B(a[14]), .C(n342), .Z(n340) );
  GTECH_XNOR2 U184 ( .A(a[15]), .B(b[15]), .Z(n337) );
  GTECH_AO21 U185 ( .A(n343), .B(n341), .C(n344), .Z(sum[14]) );
  GTECH_NOT U186 ( .A(n345), .Z(n344) );
  GTECH_MUX2 U187 ( .A(n346), .B(n347), .S(b[14]), .Z(n345) );
  GTECH_OR2 U188 ( .A(a[14]), .B(n343), .Z(n347) );
  GTECH_XNOR2 U189 ( .A(a[14]), .B(n343), .Z(n346) );
  GTECH_AO21 U190 ( .A(n348), .B(n336), .C(n342), .Z(n343) );
  GTECH_AO22 U191 ( .A(a[13]), .B(b[13]), .C(n349), .D(n350), .Z(n342) );
  GTECH_NOT U192 ( .A(n351), .Z(n349) );
  GTECH_MUX2 U193 ( .A(n352), .B(n353), .S(n336), .Z(sum[13]) );
  GTECH_XOR2 U194 ( .A(n354), .B(n355), .Z(n353) );
  GTECH_NOT U195 ( .A(n356), .Z(n354) );
  GTECH_XOR2 U196 ( .A(n355), .B(n350), .Z(n352) );
  GTECH_AOI21 U197 ( .A(a[13]), .B(b[13]), .C(n351), .Z(n355) );
  GTECH_XNOR2 U198 ( .A(n357), .B(n336), .Z(sum[12]) );
  GTECH_MUX2 U199 ( .A(n358), .B(n359), .S(n279), .Z(sum[11]) );
  GTECH_NOT U200 ( .A(n360), .Z(n279) );
  GTECH_XNOR2 U201 ( .A(n361), .B(n362), .Z(n359) );
  GTECH_AND2 U202 ( .A(n363), .B(n364), .Z(n362) );
  GTECH_OAI21 U203 ( .A(b[10]), .B(a[10]), .C(n365), .Z(n363) );
  GTECH_XOR2 U204 ( .A(n361), .B(n366), .Z(n358) );
  GTECH_XOR2 U205 ( .A(a[11]), .B(b[11]), .Z(n361) );
  GTECH_OAI21 U206 ( .A(n367), .B(n364), .C(n368), .Z(sum[10]) );
  GTECH_MUX2 U207 ( .A(n369), .B(n370), .S(b[10]), .Z(n368) );
  GTECH_OR_NOT U208 ( .A(a[10]), .B(n367), .Z(n370) );
  GTECH_XOR2 U209 ( .A(a[10]), .B(n367), .Z(n369) );
  GTECH_NOT U210 ( .A(n371), .Z(n364) );
  GTECH_AOI21 U211 ( .A(n372), .B(n360), .C(n365), .Z(n367) );
  GTECH_OAI2N2 U212 ( .A(n283), .B(n281), .C(a[9]), .D(b[9]), .Z(n365) );
  GTECH_XOR2 U213 ( .A(cin), .B(n373), .Z(sum[0]) );
  GTECH_NOT U214 ( .A(n374), .Z(cout) );
  GTECH_MUX2 U215 ( .A(n357), .B(n375), .S(n336), .Z(n374) );
  GTECH_MUX2 U216 ( .A(n284), .B(n376), .S(n360), .Z(n336) );
  GTECH_MUX2 U217 ( .A(n377), .B(n312), .S(n287), .Z(n360) );
  GTECH_NOT U218 ( .A(n301), .Z(n287) );
  GTECH_MUX2 U219 ( .A(n373), .B(n378), .S(cin), .Z(n301) );
  GTECH_OA21 U220 ( .A(a[3]), .B(n316), .C(n379), .Z(n378) );
  GTECH_AO21 U221 ( .A(n316), .B(a[3]), .C(b[3]), .Z(n379) );
  GTECH_AO21 U222 ( .A(n323), .B(a[2]), .C(n380), .Z(n316) );
  GTECH_OA21 U223 ( .A(a[2]), .B(n323), .C(b[2]), .Z(n380) );
  GTECH_AO21 U224 ( .A(n324), .B(n333), .C(n326), .Z(n323) );
  GTECH_AND2 U225 ( .A(a[1]), .B(b[1]), .Z(n326) );
  GTECH_OR2 U226 ( .A(b[1]), .B(a[1]), .Z(n324) );
  GTECH_AND2 U227 ( .A(n333), .B(n331), .Z(n373) );
  GTECH_NOT U228 ( .A(n325), .Z(n331) );
  GTECH_AND2 U229 ( .A(a[0]), .B(b[0]), .Z(n325) );
  GTECH_NOT U230 ( .A(n332), .Z(n333) );
  GTECH_NOR2 U231 ( .A(a[0]), .B(b[0]), .Z(n332) );
  GTECH_XOR2 U232 ( .A(n302), .B(n306), .Z(n312) );
  GTECH_OA21 U233 ( .A(a[7]), .B(n293), .C(n381), .Z(n377) );
  GTECH_AO21 U234 ( .A(n293), .B(a[7]), .C(b[7]), .Z(n381) );
  GTECH_AO21 U235 ( .A(n300), .B(n382), .C(n291), .Z(n293) );
  GTECH_AND2 U236 ( .A(b[6]), .B(a[6]), .Z(n291) );
  GTECH_OR_NOT U237 ( .A(b[6]), .B(n299), .Z(n382) );
  GTECH_NOT U238 ( .A(a[6]), .Z(n299) );
  GTECH_OAI21 U239 ( .A(n305), .B(n311), .C(n304), .Z(n300) );
  GTECH_OR_NOT U240 ( .A(n383), .B(b[5]), .Z(n304) );
  GTECH_NOT U241 ( .A(a[5]), .Z(n383) );
  GTECH_AND2 U242 ( .A(n302), .B(n306), .Z(n311) );
  GTECH_NOT U243 ( .A(b[4]), .Z(n306) );
  GTECH_NOT U244 ( .A(a[4]), .Z(n302) );
  GTECH_NOR2 U245 ( .A(a[5]), .B(b[5]), .Z(n305) );
  GTECH_AO21 U246 ( .A(n366), .B(a[11]), .C(n384), .Z(n376) );
  GTECH_OA21 U247 ( .A(a[11]), .B(n366), .C(b[11]), .Z(n384) );
  GTECH_AO21 U248 ( .A(n372), .B(n385), .C(n371), .Z(n366) );
  GTECH_AND2 U249 ( .A(b[10]), .B(a[10]), .Z(n371) );
  GTECH_OR2 U250 ( .A(b[10]), .B(a[10]), .Z(n385) );
  GTECH_OAI2N2 U251 ( .A(n282), .B(n283), .C(a[9]), .D(b[9]), .Z(n372) );
  GTECH_NOR2 U252 ( .A(b[9]), .B(a[9]), .Z(n283) );
  GTECH_AND_NOT U253 ( .A(n281), .B(n282), .Z(n284) );
  GTECH_AND_NOT U254 ( .A(n386), .B(b[8]), .Z(n282) );
  GTECH_OR_NOT U255 ( .A(n386), .B(b[8]), .Z(n281) );
  GTECH_NOT U256 ( .A(a[8]), .Z(n386) );
  GTECH_AOI21 U257 ( .A(n338), .B(a[15]), .C(n387), .Z(n375) );
  GTECH_OA21 U258 ( .A(a[15]), .B(n338), .C(b[15]), .Z(n387) );
  GTECH_AO21 U259 ( .A(n348), .B(n388), .C(n341), .Z(n338) );
  GTECH_AND2 U260 ( .A(b[14]), .B(a[14]), .Z(n341) );
  GTECH_OR2 U261 ( .A(b[14]), .B(a[14]), .Z(n388) );
  GTECH_OAI2N2 U262 ( .A(n356), .B(n351), .C(a[13]), .D(b[13]), .Z(n348) );
  GTECH_NOR2 U263 ( .A(a[13]), .B(b[13]), .Z(n351) );
  GTECH_OR2 U264 ( .A(n350), .B(n356), .Z(n357) );
  GTECH_NOR2 U265 ( .A(b[12]), .B(a[12]), .Z(n356) );
  GTECH_AND2 U266 ( .A(a[12]), .B(b[12]), .Z(n350) );
endmodule

