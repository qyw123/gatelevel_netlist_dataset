
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378;

  GTECH_MUX2 U130 ( .A(n269), .B(n270), .S(n271), .Z(sum[9]) );
  GTECH_XOR2 U131 ( .A(n272), .B(n273), .Z(n270) );
  GTECH_XOR2 U132 ( .A(n274), .B(n273), .Z(n269) );
  GTECH_OA21 U133 ( .A(a[9]), .B(b[9]), .C(n275), .Z(n273) );
  GTECH_OAI21 U134 ( .A(n276), .B(n277), .C(n278), .Z(sum[8]) );
  GTECH_NOT U135 ( .A(n279), .Z(n278) );
  GTECH_MUX2 U136 ( .A(n280), .B(n281), .S(n282), .Z(sum[7]) );
  GTECH_XOR2 U137 ( .A(n283), .B(n284), .Z(n281) );
  GTECH_OA21 U138 ( .A(a[6]), .B(n285), .C(n286), .Z(n283) );
  GTECH_NOT U139 ( .A(n287), .Z(n286) );
  GTECH_AOI21 U140 ( .A(n285), .B(a[6]), .C(b[6]), .Z(n287) );
  GTECH_XOR2 U141 ( .A(n284), .B(n288), .Z(n280) );
  GTECH_XNOR2 U142 ( .A(n289), .B(b[7]), .Z(n284) );
  GTECH_MUX2 U143 ( .A(n290), .B(n291), .S(n282), .Z(sum[6]) );
  GTECH_XNOR2 U144 ( .A(n292), .B(n285), .Z(n291) );
  GTECH_OAI21 U145 ( .A(n293), .B(n294), .C(n295), .Z(n285) );
  GTECH_XNOR2 U146 ( .A(n292), .B(n296), .Z(n290) );
  GTECH_XNOR2 U147 ( .A(a[6]), .B(b[6]), .Z(n292) );
  GTECH_NOT U148 ( .A(n297), .Z(sum[5]) );
  GTECH_MUX2 U149 ( .A(n298), .B(n299), .S(n300), .Z(n297) );
  GTECH_AND_NOT U150 ( .A(n295), .B(n293), .Z(n300) );
  GTECH_ADD_ABC U151 ( .A(a[4]), .B(n301), .C(b[4]), .COUT(n299) );
  GTECH_MUX2 U152 ( .A(n302), .B(n303), .S(n304), .Z(n301) );
  GTECH_OAI21 U153 ( .A(n305), .B(n306), .C(n307), .Z(n302) );
  GTECH_OA21 U154 ( .A(n308), .B(n282), .C(n294), .Z(n298) );
  GTECH_NAND2 U155 ( .A(b[4]), .B(a[4]), .Z(n294) );
  GTECH_XNOR2 U156 ( .A(n282), .B(n309), .Z(sum[4]) );
  GTECH_MUX2 U157 ( .A(n310), .B(n311), .S(n304), .Z(sum[3]) );
  GTECH_XOR2 U158 ( .A(n312), .B(n313), .Z(n311) );
  GTECH_OA21 U159 ( .A(a[2]), .B(n314), .C(n315), .Z(n312) );
  GTECH_NOT U160 ( .A(n316), .Z(n315) );
  GTECH_AOI21 U161 ( .A(n314), .B(a[2]), .C(b[2]), .Z(n316) );
  GTECH_XNOR2 U162 ( .A(n313), .B(n305), .Z(n310) );
  GTECH_XOR2 U163 ( .A(a[3]), .B(b[3]), .Z(n313) );
  GTECH_MUX2 U164 ( .A(n317), .B(n318), .S(n304), .Z(sum[2]) );
  GTECH_XNOR2 U165 ( .A(n319), .B(n314), .Z(n318) );
  GTECH_OAI21 U166 ( .A(n320), .B(n321), .C(n322), .Z(n314) );
  GTECH_XNOR2 U167 ( .A(n319), .B(n323), .Z(n317) );
  GTECH_XNOR2 U168 ( .A(a[2]), .B(b[2]), .Z(n319) );
  GTECH_MUX2 U169 ( .A(n324), .B(n325), .S(n326), .Z(sum[1]) );
  GTECH_AND_NOT U170 ( .A(n322), .B(n320), .Z(n326) );
  GTECH_NOT U171 ( .A(n327), .Z(n325) );
  GTECH_AOI21 U172 ( .A(n304), .B(n321), .C(n328), .Z(n327) );
  GTECH_OAI21 U173 ( .A(n328), .B(n304), .C(n321), .Z(n324) );
  GTECH_MUX2 U174 ( .A(n329), .B(n330), .S(n331), .Z(sum[15]) );
  GTECH_XNOR2 U175 ( .A(n332), .B(n333), .Z(n330) );
  GTECH_XNOR2 U176 ( .A(n334), .B(n332), .Z(n329) );
  GTECH_XNOR2 U177 ( .A(a[15]), .B(b[15]), .Z(n332) );
  GTECH_ADD_ABC U178 ( .A(a[14]), .B(n335), .C(b[14]), .COUT(n334) );
  GTECH_MUX2 U179 ( .A(n336), .B(n337), .S(n331), .Z(sum[14]) );
  GTECH_XOR2 U180 ( .A(n338), .B(n339), .Z(n337) );
  GTECH_XOR2 U181 ( .A(n335), .B(n339), .Z(n336) );
  GTECH_XOR2 U182 ( .A(a[14]), .B(b[14]), .Z(n339) );
  GTECH_OA21 U183 ( .A(n340), .B(n341), .C(n342), .Z(n335) );
  GTECH_MUX2 U184 ( .A(n343), .B(n344), .S(n331), .Z(sum[13]) );
  GTECH_XOR2 U185 ( .A(n345), .B(n346), .Z(n344) );
  GTECH_XOR2 U186 ( .A(n341), .B(n346), .Z(n343) );
  GTECH_AOI21 U187 ( .A(n347), .B(n348), .C(n340), .Z(n346) );
  GTECH_NAND2 U188 ( .A(n349), .B(n350), .Z(sum[12]) );
  GTECH_OAI21 U189 ( .A(n341), .B(n351), .C(n331), .Z(n349) );
  GTECH_MUX2 U190 ( .A(n352), .B(n353), .S(n271), .Z(sum[11]) );
  GTECH_XNOR2 U191 ( .A(n354), .B(n355), .Z(n353) );
  GTECH_XNOR2 U192 ( .A(n356), .B(n354), .Z(n352) );
  GTECH_XNOR2 U193 ( .A(a[11]), .B(b[11]), .Z(n354) );
  GTECH_ADD_ABC U194 ( .A(a[10]), .B(n357), .C(b[10]), .COUT(n356) );
  GTECH_MUX2 U195 ( .A(n358), .B(n359), .S(n271), .Z(sum[10]) );
  GTECH_XOR2 U196 ( .A(n360), .B(n361), .Z(n359) );
  GTECH_XOR2 U197 ( .A(n357), .B(n361), .Z(n358) );
  GTECH_XOR2 U198 ( .A(a[10]), .B(b[10]), .Z(n361) );
  GTECH_OA21 U199 ( .A(n362), .B(n274), .C(n363), .Z(n357) );
  GTECH_NOT U200 ( .A(n364), .Z(n274) );
  GTECH_XNOR2 U201 ( .A(n304), .B(n303), .Z(sum[0]) );
  GTECH_NOT U202 ( .A(n365), .Z(n303) );
  GTECH_OAI21 U203 ( .A(n366), .B(n367), .C(n350), .Z(cout) );
  GTECH_OR3 U204 ( .A(n341), .B(n351), .C(n331), .Z(n350) );
  GTECH_NOT U205 ( .A(n366), .Z(n331) );
  GTECH_AND2 U206 ( .A(a[12]), .B(b[12]), .Z(n341) );
  GTECH_AOI21 U207 ( .A(n333), .B(a[15]), .C(n368), .Z(n367) );
  GTECH_OA21 U208 ( .A(a[15]), .B(n333), .C(b[15]), .Z(n368) );
  GTECH_ADD_ABC U209 ( .A(a[14]), .B(n338), .C(b[14]), .COUT(n333) );
  GTECH_OA21 U210 ( .A(n340), .B(n345), .C(n342), .Z(n338) );
  GTECH_OR_NOT U211 ( .A(a[13]), .B(n348), .Z(n342) );
  GTECH_NOT U212 ( .A(b[13]), .Z(n348) );
  GTECH_NOT U213 ( .A(n351), .Z(n345) );
  GTECH_NOR2 U214 ( .A(a[12]), .B(b[12]), .Z(n351) );
  GTECH_AND_NOT U215 ( .A(b[13]), .B(n347), .Z(n340) );
  GTECH_NOT U216 ( .A(a[13]), .Z(n347) );
  GTECH_AOI21 U217 ( .A(n271), .B(n369), .C(n279), .Z(n366) );
  GTECH_AND2 U218 ( .A(n276), .B(n277), .Z(n279) );
  GTECH_NOT U219 ( .A(n271), .Z(n277) );
  GTECH_AND2 U220 ( .A(n272), .B(n364), .Z(n276) );
  GTECH_NAND2 U221 ( .A(a[8]), .B(b[8]), .Z(n364) );
  GTECH_OA21 U222 ( .A(a[11]), .B(n355), .C(n370), .Z(n369) );
  GTECH_NOT U223 ( .A(n371), .Z(n370) );
  GTECH_AOI21 U224 ( .A(n355), .B(a[11]), .C(b[11]), .Z(n371) );
  GTECH_ADD_ABC U225 ( .A(n360), .B(a[10]), .C(b[10]), .COUT(n355) );
  GTECH_OA21 U226 ( .A(n362), .B(n272), .C(n363), .Z(n360) );
  GTECH_OR2 U227 ( .A(a[9]), .B(b[9]), .Z(n363) );
  GTECH_OR2 U228 ( .A(a[8]), .B(b[8]), .Z(n272) );
  GTECH_NOT U229 ( .A(n275), .Z(n362) );
  GTECH_NAND2 U230 ( .A(b[9]), .B(a[9]), .Z(n275) );
  GTECH_MUX2 U231 ( .A(n372), .B(n309), .S(n282), .Z(n271) );
  GTECH_MUX2 U232 ( .A(n373), .B(n365), .S(n304), .Z(n282) );
  GTECH_NOT U233 ( .A(cin), .Z(n304) );
  GTECH_OR_NOT U234 ( .A(n328), .B(n321), .Z(n365) );
  GTECH_NAND2 U235 ( .A(b[0]), .B(a[0]), .Z(n321) );
  GTECH_OA21 U236 ( .A(n305), .B(n306), .C(n307), .Z(n373) );
  GTECH_OAI21 U237 ( .A(a[3]), .B(n374), .C(b[3]), .Z(n307) );
  GTECH_NOT U238 ( .A(n305), .Z(n374) );
  GTECH_NOT U239 ( .A(a[3]), .Z(n306) );
  GTECH_AOI21 U240 ( .A(n323), .B(a[2]), .C(n375), .Z(n305) );
  GTECH_OA21 U241 ( .A(a[2]), .B(n323), .C(b[2]), .Z(n375) );
  GTECH_OAI21 U242 ( .A(n328), .B(n320), .C(n322), .Z(n323) );
  GTECH_NAND2 U243 ( .A(a[1]), .B(b[1]), .Z(n322) );
  GTECH_NOR2 U244 ( .A(b[1]), .B(a[1]), .Z(n320) );
  GTECH_NOR2 U245 ( .A(a[0]), .B(b[0]), .Z(n328) );
  GTECH_XOR2 U246 ( .A(a[4]), .B(b[4]), .Z(n309) );
  GTECH_AOI21 U247 ( .A(n289), .B(n376), .C(n377), .Z(n372) );
  GTECH_AOI21 U248 ( .A(n288), .B(a[7]), .C(b[7]), .Z(n377) );
  GTECH_NOT U249 ( .A(n376), .Z(n288) );
  GTECH_AOI21 U250 ( .A(n296), .B(a[6]), .C(n378), .Z(n376) );
  GTECH_OA21 U251 ( .A(a[6]), .B(n296), .C(b[6]), .Z(n378) );
  GTECH_OAI21 U252 ( .A(n308), .B(n293), .C(n295), .Z(n296) );
  GTECH_NAND2 U253 ( .A(b[5]), .B(a[5]), .Z(n295) );
  GTECH_NOR2 U254 ( .A(b[5]), .B(a[5]), .Z(n293) );
  GTECH_NOR2 U255 ( .A(b[4]), .B(a[4]), .Z(n308) );
  GTECH_NOT U256 ( .A(a[7]), .Z(n289) );
endmodule

