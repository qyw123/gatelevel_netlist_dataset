
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373;

  GTECH_MUX2 U136 ( .A(n275), .B(n276), .S(n277), .Z(sum[9]) );
  GTECH_XOR2 U137 ( .A(n278), .B(n279), .Z(n276) );
  GTECH_XOR2 U138 ( .A(n279), .B(n280), .Z(n275) );
  GTECH_OA21 U139 ( .A(a[9]), .B(b[9]), .C(n281), .Z(n279) );
  GTECH_OAI21 U140 ( .A(n282), .B(n283), .C(n284), .Z(sum[8]) );
  GTECH_MUX2 U141 ( .A(n285), .B(n286), .S(n287), .Z(sum[7]) );
  GTECH_XOR2 U142 ( .A(n288), .B(n289), .Z(n286) );
  GTECH_OA21 U143 ( .A(n290), .B(n291), .C(n292), .Z(n289) );
  GTECH_XNOR2 U144 ( .A(n288), .B(n293), .Z(n285) );
  GTECH_XNOR2 U145 ( .A(a[7]), .B(b[7]), .Z(n288) );
  GTECH_MUX2 U146 ( .A(n294), .B(n295), .S(n287), .Z(sum[6]) );
  GTECH_XNOR2 U147 ( .A(n296), .B(n291), .Z(n295) );
  GTECH_OA21 U148 ( .A(n297), .B(n298), .C(n299), .Z(n291) );
  GTECH_XNOR2 U149 ( .A(n296), .B(n300), .Z(n294) );
  GTECH_AND_NOT U150 ( .A(n292), .B(n290), .Z(n296) );
  GTECH_MUX2 U151 ( .A(n301), .B(n302), .S(n303), .Z(sum[5]) );
  GTECH_AND_NOT U152 ( .A(n299), .B(n297), .Z(n303) );
  GTECH_AO21 U153 ( .A(n298), .B(n287), .C(n304), .Z(n302) );
  GTECH_OAI21 U154 ( .A(n304), .B(n287), .C(n298), .Z(n301) );
  GTECH_XNOR2 U155 ( .A(n305), .B(n287), .Z(sum[4]) );
  GTECH_MUX2 U156 ( .A(n306), .B(n307), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U157 ( .A(n308), .B(n309), .Z(n307) );
  GTECH_XOR2 U158 ( .A(n308), .B(n310), .Z(n306) );
  GTECH_OA21 U159 ( .A(n311), .B(n312), .C(n313), .Z(n310) );
  GTECH_XNOR2 U160 ( .A(a[3]), .B(b[3]), .Z(n308) );
  GTECH_MUX2 U161 ( .A(n314), .B(n315), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U162 ( .A(n316), .B(n317), .Z(n315) );
  GTECH_XNOR2 U163 ( .A(n312), .B(n316), .Z(n314) );
  GTECH_AND_NOT U164 ( .A(n313), .B(n311), .Z(n316) );
  GTECH_AOI21 U165 ( .A(n318), .B(n319), .C(n320), .Z(n312) );
  GTECH_MUX2 U166 ( .A(n321), .B(n322), .S(n323), .Z(sum[1]) );
  GTECH_AND_NOT U167 ( .A(n318), .B(n320), .Z(n323) );
  GTECH_OAI21 U168 ( .A(cin), .B(n319), .C(n324), .Z(n322) );
  GTECH_AO21 U169 ( .A(n324), .B(cin), .C(n319), .Z(n321) );
  GTECH_MUX2 U170 ( .A(n325), .B(n326), .S(n327), .Z(sum[15]) );
  GTECH_XOR2 U171 ( .A(n328), .B(n329), .Z(n326) );
  GTECH_XOR2 U172 ( .A(n330), .B(n329), .Z(n325) );
  GTECH_XOR2 U173 ( .A(a[15]), .B(b[15]), .Z(n329) );
  GTECH_OA21 U174 ( .A(n331), .B(n332), .C(n333), .Z(n330) );
  GTECH_MUX2 U175 ( .A(n334), .B(n335), .S(n327), .Z(sum[14]) );
  GTECH_XNOR2 U176 ( .A(n336), .B(n337), .Z(n335) );
  GTECH_XNOR2 U177 ( .A(n336), .B(n332), .Z(n334) );
  GTECH_AOI21 U178 ( .A(n338), .B(n339), .C(n340), .Z(n332) );
  GTECH_OAI21 U179 ( .A(a[14]), .B(b[14]), .C(n341), .Z(n336) );
  GTECH_MUX2 U180 ( .A(n342), .B(n343), .S(n327), .Z(sum[13]) );
  GTECH_XOR2 U181 ( .A(n344), .B(n345), .Z(n343) );
  GTECH_XOR2 U182 ( .A(n345), .B(n339), .Z(n342) );
  GTECH_NOT U183 ( .A(n346), .Z(n339) );
  GTECH_OAI21 U184 ( .A(a[13]), .B(b[13]), .C(n338), .Z(n345) );
  GTECH_NAND2 U185 ( .A(n347), .B(n348), .Z(sum[12]) );
  GTECH_OAI21 U186 ( .A(n346), .B(n344), .C(n327), .Z(n347) );
  GTECH_MUX2 U187 ( .A(n349), .B(n350), .S(n277), .Z(sum[11]) );
  GTECH_XNOR2 U188 ( .A(n351), .B(n352), .Z(n350) );
  GTECH_XOR2 U189 ( .A(n351), .B(n353), .Z(n349) );
  GTECH_AOI21 U190 ( .A(n354), .B(n355), .C(n356), .Z(n353) );
  GTECH_XNOR2 U191 ( .A(a[11]), .B(b[11]), .Z(n351) );
  GTECH_MUX2 U192 ( .A(n357), .B(n358), .S(n277), .Z(sum[10]) );
  GTECH_XOR2 U193 ( .A(n359), .B(n360), .Z(n358) );
  GTECH_XOR2 U194 ( .A(n359), .B(n355), .Z(n357) );
  GTECH_OA21 U195 ( .A(n361), .B(n280), .C(n362), .Z(n355) );
  GTECH_AND_NOT U196 ( .A(n354), .B(n356), .Z(n359) );
  GTECH_XNOR2 U197 ( .A(cin), .B(n363), .Z(sum[0]) );
  GTECH_OAI21 U198 ( .A(n364), .B(n365), .C(n348), .Z(cout) );
  GTECH_OR3 U199 ( .A(n344), .B(n346), .C(n327), .Z(n348) );
  GTECH_NOT U200 ( .A(n364), .Z(n327) );
  GTECH_AND2 U201 ( .A(b[12]), .B(a[12]), .Z(n346) );
  GTECH_AOI21 U202 ( .A(a[15]), .B(n328), .C(n366), .Z(n365) );
  GTECH_OA21 U203 ( .A(n328), .B(a[15]), .C(b[15]), .Z(n366) );
  GTECH_OA21 U204 ( .A(n331), .B(n337), .C(n333), .Z(n328) );
  GTECH_OR2 U205 ( .A(b[14]), .B(a[14]), .Z(n333) );
  GTECH_AOI21 U206 ( .A(n338), .B(n344), .C(n340), .Z(n337) );
  GTECH_NOR2 U207 ( .A(b[13]), .B(a[13]), .Z(n340) );
  GTECH_NOR2 U208 ( .A(a[12]), .B(b[12]), .Z(n344) );
  GTECH_NAND2 U209 ( .A(a[13]), .B(b[13]), .Z(n338) );
  GTECH_NOT U210 ( .A(n341), .Z(n331) );
  GTECH_NAND2 U211 ( .A(a[14]), .B(b[14]), .Z(n341) );
  GTECH_OA21 U212 ( .A(n283), .B(n367), .C(n284), .Z(n364) );
  GTECH_NAND2 U213 ( .A(n283), .B(n282), .Z(n284) );
  GTECH_AND_NOT U214 ( .A(n278), .B(n280), .Z(n282) );
  GTECH_AND2 U215 ( .A(b[8]), .B(a[8]), .Z(n280) );
  GTECH_OAI21 U216 ( .A(a[11]), .B(n352), .C(n368), .Z(n367) );
  GTECH_AO21 U217 ( .A(n352), .B(a[11]), .C(b[11]), .Z(n368) );
  GTECH_AO21 U218 ( .A(n354), .B(n360), .C(n356), .Z(n352) );
  GTECH_AND2 U219 ( .A(a[10]), .B(b[10]), .Z(n356) );
  GTECH_OA21 U220 ( .A(n361), .B(n278), .C(n362), .Z(n360) );
  GTECH_OR2 U221 ( .A(b[9]), .B(a[9]), .Z(n362) );
  GTECH_OR2 U222 ( .A(a[8]), .B(b[8]), .Z(n278) );
  GTECH_NOT U223 ( .A(n281), .Z(n361) );
  GTECH_NAND2 U224 ( .A(b[9]), .B(a[9]), .Z(n281) );
  GTECH_OR2 U225 ( .A(a[10]), .B(b[10]), .Z(n354) );
  GTECH_NOT U226 ( .A(n277), .Z(n283) );
  GTECH_MUX2 U227 ( .A(n369), .B(n305), .S(n287), .Z(n277) );
  GTECH_MUX2 U228 ( .A(n363), .B(n370), .S(cin), .Z(n287) );
  GTECH_AOI21 U229 ( .A(n309), .B(a[3]), .C(n371), .Z(n370) );
  GTECH_OA21 U230 ( .A(a[3]), .B(n309), .C(b[3]), .Z(n371) );
  GTECH_OAI21 U231 ( .A(n317), .B(n311), .C(n313), .Z(n309) );
  GTECH_NAND2 U232 ( .A(b[2]), .B(a[2]), .Z(n313) );
  GTECH_NOR2 U233 ( .A(a[2]), .B(b[2]), .Z(n311) );
  GTECH_AOI21 U234 ( .A(n318), .B(n324), .C(n320), .Z(n317) );
  GTECH_AND2 U235 ( .A(b[1]), .B(a[1]), .Z(n320) );
  GTECH_OR2 U236 ( .A(b[1]), .B(a[1]), .Z(n318) );
  GTECH_NAND2 U237 ( .A(n324), .B(n372), .Z(n363) );
  GTECH_NOT U238 ( .A(n319), .Z(n372) );
  GTECH_AND2 U239 ( .A(b[0]), .B(a[0]), .Z(n319) );
  GTECH_OR2 U240 ( .A(a[0]), .B(b[0]), .Z(n324) );
  GTECH_AND_NOT U241 ( .A(n298), .B(n304), .Z(n305) );
  GTECH_NAND2 U242 ( .A(b[4]), .B(a[4]), .Z(n298) );
  GTECH_OA21 U243 ( .A(a[7]), .B(n293), .C(n373), .Z(n369) );
  GTECH_AO21 U244 ( .A(n293), .B(a[7]), .C(b[7]), .Z(n373) );
  GTECH_OAI21 U245 ( .A(n300), .B(n290), .C(n292), .Z(n293) );
  GTECH_NAND2 U246 ( .A(b[6]), .B(a[6]), .Z(n292) );
  GTECH_NOR2 U247 ( .A(a[6]), .B(b[6]), .Z(n290) );
  GTECH_OA21 U248 ( .A(n304), .B(n297), .C(n299), .Z(n300) );
  GTECH_NAND2 U249 ( .A(b[5]), .B(a[5]), .Z(n299) );
  GTECH_NOR2 U250 ( .A(b[5]), .B(a[5]), .Z(n297) );
  GTECH_NOR2 U251 ( .A(b[4]), .B(a[4]), .Z(n304) );
endmodule

