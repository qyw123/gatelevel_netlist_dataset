
module carry_select_adder8 ( a, b, cin, cout, sum );
  input [7:0] a;
  input [7:0] b;
  output [7:0] sum;
  input cin;
  output cout;
  wire   n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189;

  GTECH_MUX2 U64 ( .A(n133), .B(n134), .S(n135), .Z(sum[7]) );
  GTECH_XNOR2 U65 ( .A(n136), .B(n137), .Z(n134) );
  GTECH_XNOR2 U66 ( .A(n136), .B(n138), .Z(n133) );
  GTECH_AOI21 U67 ( .A(n139), .B(n140), .C(n141), .Z(n138) );
  GTECH_NOT U68 ( .A(n142), .Z(n141) );
  GTECH_OR2 U69 ( .A(a[6]), .B(b[6]), .Z(n139) );
  GTECH_XNOR2 U70 ( .A(a[7]), .B(n143), .Z(n136) );
  GTECH_MUX2 U71 ( .A(n144), .B(n145), .S(n135), .Z(sum[6]) );
  GTECH_XOR2 U72 ( .A(n146), .B(n147), .Z(n145) );
  GTECH_XOR2 U73 ( .A(n146), .B(n140), .Z(n144) );
  GTECH_OR_NOT U74 ( .A(n148), .B(n149), .Z(n140) );
  GTECH_OAI21 U75 ( .A(b[5]), .B(a[5]), .C(n150), .Z(n149) );
  GTECH_OA21 U76 ( .A(b[6]), .B(a[6]), .C(n142), .Z(n146) );
  GTECH_MUX2 U77 ( .A(n151), .B(n152), .S(n135), .Z(sum[5]) );
  GTECH_XOR2 U78 ( .A(n153), .B(n154), .Z(n152) );
  GTECH_XNOR2 U79 ( .A(n150), .B(n153), .Z(n151) );
  GTECH_AO21 U80 ( .A(n155), .B(n156), .C(n148), .Z(n153) );
  GTECH_NAND2 U81 ( .A(n157), .B(n158), .Z(sum[4]) );
  GTECH_OAI21 U82 ( .A(n150), .B(n154), .C(n135), .Z(n158) );
  GTECH_MUX2 U83 ( .A(n159), .B(n160), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U84 ( .A(n161), .B(n162), .Z(n160) );
  GTECH_XNOR2 U85 ( .A(n161), .B(n163), .Z(n159) );
  GTECH_AOI21 U86 ( .A(n164), .B(n165), .C(n166), .Z(n163) );
  GTECH_NOT U87 ( .A(n167), .Z(n166) );
  GTECH_OR2 U88 ( .A(a[2]), .B(b[2]), .Z(n164) );
  GTECH_XOR2 U89 ( .A(a[3]), .B(b[3]), .Z(n161) );
  GTECH_MUX2 U90 ( .A(n168), .B(n169), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U91 ( .A(n170), .B(n171), .Z(n169) );
  GTECH_XOR2 U92 ( .A(n170), .B(n165), .Z(n168) );
  GTECH_NAND2 U93 ( .A(n172), .B(n173), .Z(n165) );
  GTECH_OAI21 U94 ( .A(b[1]), .B(a[1]), .C(n174), .Z(n173) );
  GTECH_OA21 U95 ( .A(b[2]), .B(a[2]), .C(n167), .Z(n170) );
  GTECH_MUX2 U96 ( .A(n175), .B(n176), .S(n177), .Z(sum[1]) );
  GTECH_OA21 U97 ( .A(b[1]), .B(a[1]), .C(n172), .Z(n177) );
  GTECH_OAI21 U98 ( .A(cin), .B(n174), .C(n178), .Z(n176) );
  GTECH_AO21 U99 ( .A(n178), .B(cin), .C(n174), .Z(n175) );
  GTECH_ADD_AB U100 ( .A(a[0]), .B(b[0]), .COUT(n174) );
  GTECH_XOR2 U101 ( .A(cin), .B(n179), .Z(sum[0]) );
  GTECH_OAI21 U102 ( .A(n180), .B(n181), .C(n157), .Z(cout) );
  GTECH_OR3 U103 ( .A(n150), .B(n154), .C(n135), .Z(n157) );
  GTECH_ADD_AB U104 ( .A(b[4]), .B(a[4]), .COUT(n150) );
  GTECH_NOT U105 ( .A(n135), .Z(n181) );
  GTECH_MUX2 U106 ( .A(n179), .B(n182), .S(cin), .Z(n135) );
  GTECH_OA21 U107 ( .A(a[3]), .B(n162), .C(n183), .Z(n182) );
  GTECH_AO21 U108 ( .A(n162), .B(a[3]), .C(b[3]), .Z(n183) );
  GTECH_NAND2 U109 ( .A(n167), .B(n184), .Z(n162) );
  GTECH_OAI21 U110 ( .A(a[2]), .B(b[2]), .C(n171), .Z(n184) );
  GTECH_NAND2 U111 ( .A(n172), .B(n185), .Z(n171) );
  GTECH_OAI21 U112 ( .A(a[1]), .B(b[1]), .C(n178), .Z(n185) );
  GTECH_OR2 U113 ( .A(a[0]), .B(b[0]), .Z(n178) );
  GTECH_NAND2 U114 ( .A(b[1]), .B(a[1]), .Z(n172) );
  GTECH_NAND2 U115 ( .A(b[2]), .B(a[2]), .Z(n167) );
  GTECH_XOR2 U116 ( .A(a[0]), .B(b[0]), .Z(n179) );
  GTECH_OA21 U117 ( .A(n137), .B(n186), .C(n187), .Z(n180) );
  GTECH_AO21 U118 ( .A(n186), .B(n137), .C(n143), .Z(n187) );
  GTECH_NOT U119 ( .A(b[7]), .Z(n143) );
  GTECH_NOT U120 ( .A(a[7]), .Z(n186) );
  GTECH_ADD_AB U121 ( .A(n142), .B(n188), .COUT(n137) );
  GTECH_OAI21 U122 ( .A(a[6]), .B(b[6]), .C(n147), .Z(n188) );
  GTECH_OR_NOT U123 ( .A(n148), .B(n189), .Z(n147) );
  GTECH_AO21 U124 ( .A(n156), .B(n155), .C(n154), .Z(n189) );
  GTECH_NOR2 U125 ( .A(a[4]), .B(b[4]), .Z(n154) );
  GTECH_NOR2 U126 ( .A(n155), .B(n156), .Z(n148) );
  GTECH_NOT U127 ( .A(a[5]), .Z(n156) );
  GTECH_NOT U128 ( .A(b[5]), .Z(n155) );
  GTECH_NAND2 U129 ( .A(b[6]), .B(a[6]), .Z(n142) );
endmodule

