
module CRC_16_parallel ( clk, rst_n, data, data_valid, crc );
  input [7:0] data;
  output [15:0] crc;
  input clk, rst_n, data_valid;
  wire   N11, N15, N19, N23, N34, N37, N39, N41, N43, N45, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N58, N60, N62, N64, N69, N70, N99, N209,
         N222, N235, N248, N261, N274, N287, N298, N307, N316, N323, N328,
         N331, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223;
  wire   [23:0] temp;

  GTECH_FJK2S temp_reg_15_ ( .J(1'b0), .K(1'b0), .TI(N56), .TE(N287), .CP(clk), 
        .CD(rst_n), .Q(temp[15]) );
  GTECH_FJK2S temp_reg_14_ ( .J(1'b0), .K(1'b0), .TI(N55), .TE(N209), .CP(clk), 
        .CD(rst_n), .Q(temp[14]) );
  GTECH_FJK2S temp_reg_13_ ( .J(1'b0), .K(1'b0), .TI(N54), .TE(N222), .CP(clk), 
        .CD(rst_n), .Q(temp[13]) );
  GTECH_FJK2S temp_reg_12_ ( .J(1'b0), .K(1'b0), .TI(N53), .TE(N235), .CP(clk), 
        .CD(rst_n), .Q(temp[12]), .QN(N53) );
  GTECH_FJK2S temp_reg_11_ ( .J(1'b0), .K(1'b0), .TI(N52), .TE(N248), .CP(clk), 
        .CD(rst_n), .Q(temp[11]) );
  GTECH_FJK2S temp_reg_10_ ( .J(1'b0), .K(1'b0), .TI(N51), .TE(N261), .CP(clk), 
        .CD(rst_n), .Q(temp[10]) );
  GTECH_FJK2S temp_reg_9_ ( .J(1'b0), .K(1'b0), .TI(N50), .TE(N274), .CP(clk), 
        .CD(rst_n), .Q(temp[9]) );
  GTECH_FJK2S temp_reg_8_ ( .J(1'b0), .K(1'b0), .TI(N49), .TE(N287), .CP(clk), 
        .CD(rst_n), .Q(temp[8]) );
  GTECH_FJK2S temp_reg_7_ ( .J(1'b0), .K(1'b0), .TI(N48), .TE(N298), .CP(clk), 
        .CD(rst_n), .Q(temp[7]) );
  GTECH_FJK2S temp_reg_6_ ( .J(1'b0), .K(1'b0), .TI(N47), .TE(N307), .CP(clk), 
        .CD(rst_n), .Q(temp[6]) );
  GTECH_FJK2S temp_reg_5_ ( .J(1'b0), .K(1'b0), .TI(N45), .TE(N316), .CP(clk), 
        .CD(rst_n), .Q(temp[5]), .QN(N45) );
  GTECH_FJK2S temp_reg_4_ ( .J(1'b0), .K(1'b0), .TI(N43), .TE(N323), .CP(clk), 
        .CD(rst_n), .Q(temp[4]) );
  GTECH_FJK2S temp_reg_3_ ( .J(1'b0), .K(1'b0), .TI(N41), .TE(N328), .CP(clk), 
        .CD(rst_n), .Q(temp[3]) );
  GTECH_FJK2S temp_reg_2_ ( .J(1'b0), .K(1'b0), .TI(N39), .TE(N331), .CP(clk), 
        .CD(rst_n), .Q(temp[2]) );
  GTECH_FJK2S temp_reg_1_ ( .J(1'b0), .K(1'b0), .TI(N37), .TE(N70), .CP(clk), 
        .CD(rst_n), .Q(temp[1]) );
  GTECH_FJK2S temp_reg_0_ ( .J(1'b0), .K(1'b0), .TI(N34), .TE(N69), .CP(clk), 
        .CD(rst_n), .Q(temp[0]), .QN(N34) );
  GTECH_FJK2S crc_reg_15_ ( .J(1'b0), .K(1'b0), .TI(temp[15]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[15]) );
  GTECH_FJK2S crc_reg_14_ ( .J(1'b0), .K(1'b0), .TI(temp[14]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[14]) );
  GTECH_FJK2S crc_reg_13_ ( .J(1'b0), .K(1'b0), .TI(temp[13]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[13]) );
  GTECH_FJK2S crc_reg_12_ ( .J(1'b0), .K(1'b0), .TI(temp[12]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[12]) );
  GTECH_FJK2S crc_reg_11_ ( .J(1'b0), .K(1'b0), .TI(temp[11]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[11]) );
  GTECH_FJK2S crc_reg_10_ ( .J(1'b0), .K(1'b0), .TI(temp[10]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[10]) );
  GTECH_FJK2S crc_reg_9_ ( .J(1'b0), .K(1'b0), .TI(temp[9]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[9]) );
  GTECH_FJK2S crc_reg_8_ ( .J(1'b0), .K(1'b0), .TI(temp[8]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[8]) );
  GTECH_FJK2S crc_reg_7_ ( .J(1'b0), .K(1'b0), .TI(temp[7]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[7]) );
  GTECH_FJK2S crc_reg_6_ ( .J(1'b0), .K(1'b0), .TI(temp[6]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[6]) );
  GTECH_FJK2S crc_reg_5_ ( .J(1'b0), .K(1'b0), .TI(temp[5]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[5]) );
  GTECH_FJK2S crc_reg_4_ ( .J(1'b0), .K(1'b0), .TI(temp[4]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[4]) );
  GTECH_FJK2S crc_reg_3_ ( .J(1'b0), .K(1'b0), .TI(temp[3]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[3]) );
  GTECH_FJK2S crc_reg_2_ ( .J(1'b0), .K(1'b0), .TI(temp[2]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[2]) );
  GTECH_FJK2S crc_reg_1_ ( .J(1'b0), .K(1'b0), .TI(temp[1]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[1]) );
  GTECH_FJK2S crc_reg_0_ ( .J(1'b0), .K(1'b0), .TI(temp[0]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[0]) );
  GTECH_FD3 temp_reg_23_ ( .D(n99), .CP(clk), .CD(n91), .SD(n90), .Q(temp[23]), 
        .QN(N11) );
  GTECH_FD3 temp_reg_22_ ( .D(n98), .CP(clk), .CD(n89), .SD(n88), .Q(temp[22]), 
        .QN(N15) );
  GTECH_FD3 temp_reg_21_ ( .D(n97), .CP(clk), .CD(n87), .SD(n86), .Q(temp[21]), 
        .QN(N19) );
  GTECH_FD3 temp_reg_20_ ( .D(n96), .CP(clk), .CD(n85), .SD(n84), .Q(temp[20]), 
        .QN(N23) );
  GTECH_FD3 temp_reg_19_ ( .D(n95), .CP(clk), .CD(n83), .SD(n82), .Q(temp[19]), 
        .QN(N64) );
  GTECH_FD3 temp_reg_18_ ( .D(n94), .CP(clk), .CD(n81), .SD(n80), .Q(temp[18]), 
        .QN(N62) );
  GTECH_FD3 temp_reg_17_ ( .D(n93), .CP(clk), .CD(n79), .SD(n78), .Q(temp[17]), 
        .QN(N60) );
  GTECH_FD3 temp_reg_16_ ( .D(n92), .CP(clk), .CD(n77), .SD(n76), .Q(temp[16]), 
        .QN(N58) );
  GTECH_AND2 U143 ( .A(temp[23]), .B(n148), .Z(n99) );
  GTECH_OA21 U144 ( .A(temp[23]), .B(n148), .C(temp[22]), .Z(n98) );
  GTECH_AND2 U145 ( .A(temp[21]), .B(n149), .Z(n97) );
  GTECH_AND2 U146 ( .A(temp[20]), .B(n150), .Z(n96) );
  GTECH_XOR2 U147 ( .A(temp[19]), .B(n151), .Z(n95) );
  GTECH_OA21 U148 ( .A(n152), .B(temp[23]), .C(data_valid), .Z(n151) );
  GTECH_NOT U149 ( .A(n153), .Z(n152) );
  GTECH_XOR2 U150 ( .A(temp[18]), .B(n154), .Z(n94) );
  GTECH_AND3 U151 ( .A(data_valid), .B(n155), .C(n156), .Z(n154) );
  GTECH_OA21 U152 ( .A(n157), .B(temp[22]), .C(n158), .Z(n156) );
  GTECH_MUX2 U153 ( .A(n159), .B(n160), .S(temp[17]), .Z(n93) );
  GTECH_OAI21 U154 ( .A(temp[21]), .B(n161), .C(n162), .Z(n160) );
  GTECH_AND2 U155 ( .A(n162), .B(temp[21]), .Z(n159) );
  GTECH_XOR2 U156 ( .A(N274), .B(temp[16]), .Z(n92) );
  GTECH_NAND2 U157 ( .A(n163), .B(n164), .Z(n91) );
  GTECH_NOT U158 ( .A(data[7]), .Z(n164) );
  GTECH_NAND2 U159 ( .A(data[7]), .B(n163), .Z(n90) );
  GTECH_NAND2 U160 ( .A(n163), .B(n165), .Z(n89) );
  GTECH_NOT U161 ( .A(data[6]), .Z(n165) );
  GTECH_NAND2 U162 ( .A(data[6]), .B(n163), .Z(n88) );
  GTECH_NAND2 U163 ( .A(n163), .B(n166), .Z(n87) );
  GTECH_NOT U164 ( .A(data[5]), .Z(n166) );
  GTECH_NAND2 U165 ( .A(data[5]), .B(n163), .Z(n86) );
  GTECH_NAND2 U166 ( .A(n163), .B(n167), .Z(n85) );
  GTECH_NOT U167 ( .A(data[4]), .Z(n167) );
  GTECH_NAND2 U168 ( .A(data[4]), .B(n163), .Z(n84) );
  GTECH_NAND2 U169 ( .A(n163), .B(n168), .Z(n83) );
  GTECH_NOT U170 ( .A(data[3]), .Z(n168) );
  GTECH_NAND2 U171 ( .A(data[3]), .B(n163), .Z(n82) );
  GTECH_NAND2 U172 ( .A(n163), .B(n169), .Z(n81) );
  GTECH_NOT U173 ( .A(data[2]), .Z(n169) );
  GTECH_NAND2 U174 ( .A(data[2]), .B(n163), .Z(n80) );
  GTECH_NAND2 U175 ( .A(n163), .B(n170), .Z(n79) );
  GTECH_NOT U176 ( .A(data[1]), .Z(n170) );
  GTECH_NAND2 U177 ( .A(data[1]), .B(n163), .Z(n78) );
  GTECH_NAND2 U178 ( .A(n163), .B(n171), .Z(n77) );
  GTECH_NOT U179 ( .A(data[0]), .Z(n171) );
  GTECH_NAND2 U180 ( .A(data[0]), .B(n163), .Z(n76) );
  GTECH_NOT U181 ( .A(rst_n), .Z(n163) );
  GTECH_AND4 U182 ( .A(n172), .B(n173), .C(data_valid), .D(n174), .Z(N99) );
  GTECH_NOT U183 ( .A(n175), .Z(N69) );
  GTECH_XOR2 U184 ( .A(temp[19]), .B(temp[15]), .Z(N56) );
  GTECH_XOR2 U185 ( .A(temp[18]), .B(temp[14]), .Z(N55) );
  GTECH_XOR2 U186 ( .A(temp[17]), .B(temp[13]), .Z(N54) );
  GTECH_XOR2 U187 ( .A(temp[22]), .B(temp[11]), .Z(N52) );
  GTECH_XOR2 U188 ( .A(temp[21]), .B(temp[10]), .Z(N51) );
  GTECH_XOR2 U189 ( .A(temp[9]), .B(temp[20]), .Z(N50) );
  GTECH_XOR2 U190 ( .A(temp[8]), .B(temp[19]), .Z(N49) );
  GTECH_XOR2 U191 ( .A(n176), .B(temp[7]), .Z(N48) );
  GTECH_NAND2 U192 ( .A(n158), .B(n177), .Z(n176) );
  GTECH_XOR2 U193 ( .A(n178), .B(temp[6]), .Z(N47) );
  GTECH_NAND2 U194 ( .A(n179), .B(n180), .Z(n178) );
  GTECH_XOR2 U195 ( .A(temp[4]), .B(temp[20]), .Z(N43) );
  GTECH_XOR2 U196 ( .A(temp[3]), .B(temp[19]), .Z(N41) );
  GTECH_XOR2 U197 ( .A(temp[2]), .B(temp[18]), .Z(N39) );
  GTECH_XOR2 U198 ( .A(temp[1]), .B(temp[17]), .Z(N37) );
  GTECH_AND2 U199 ( .A(n181), .B(n182), .Z(N331) );
  GTECH_OA21 U200 ( .A(n172), .B(temp[19]), .C(n183), .Z(N328) );
  GTECH_AND2 U201 ( .A(n184), .B(n185), .Z(N323) );
  GTECH_OAI21 U202 ( .A(temp[19]), .B(n186), .C(n187), .Z(n185) );
  GTECH_AND2 U203 ( .A(n188), .B(n189), .Z(N316) );
  GTECH_OA21 U204 ( .A(n190), .B(n189), .C(n191), .Z(N307) );
  GTECH_OAI21 U205 ( .A(temp[21]), .B(n192), .C(n162), .Z(n191) );
  GTECH_OAI21 U206 ( .A(n157), .B(n149), .C(n193), .Z(n189) );
  GTECH_NOT U207 ( .A(n184), .Z(n193) );
  GTECH_OAI21 U208 ( .A(n187), .B(n150), .C(n194), .Z(n184) );
  GTECH_NOT U209 ( .A(n183), .Z(n194) );
  GTECH_OAI21 U210 ( .A(n148), .B(n153), .C(n195), .Z(n183) );
  GTECH_NOT U211 ( .A(n181), .Z(n195) );
  GTECH_OAI21 U212 ( .A(n148), .B(n196), .C(n197), .Z(n181) );
  GTECH_NOT U213 ( .A(N70), .Z(n197) );
  GTECH_OAI21 U214 ( .A(n148), .B(n182), .C(n175), .Z(N70) );
  GTECH_NAND2 U215 ( .A(n198), .B(data_valid), .Z(n175) );
  GTECH_NOT U216 ( .A(n199), .Z(n198) );
  GTECH_AND3 U217 ( .A(data_valid), .B(n158), .C(temp[22]), .Z(n190) );
  GTECH_OAI21 U218 ( .A(n158), .B(n148), .C(n200), .Z(N298) );
  GTECH_OR3 U219 ( .A(n201), .B(n202), .C(n203), .Z(n200) );
  GTECH_OAI22 U220 ( .A(n153), .B(n203), .C(n186), .D(n204), .Z(N287) );
  GTECH_OAI21 U221 ( .A(n187), .B(n150), .C(n205), .Z(N274) );
  GTECH_OR3 U222 ( .A(temp[19]), .B(n186), .C(n204), .Z(n205) );
  GTECH_AND3 U223 ( .A(n206), .B(n188), .C(n207), .Z(N261) );
  GTECH_OAI21 U224 ( .A(n208), .B(n186), .C(n157), .Z(n188) );
  GTECH_AND2 U225 ( .A(n209), .B(n207), .Z(N248) );
  GTECH_NOT U226 ( .A(n203), .Z(n207) );
  GTECH_OA21 U227 ( .A(n210), .B(temp[22]), .C(n158), .Z(n209) );
  GTECH_AND3 U228 ( .A(n211), .B(n157), .C(n172), .Z(n210) );
  GTECH_NOT U229 ( .A(n186), .Z(n172) );
  GTECH_OAI21 U230 ( .A(n158), .B(n148), .C(n212), .Z(N235) );
  GTECH_OR3 U231 ( .A(n202), .B(n186), .C(n203), .Z(n212) );
  GTECH_NOT U232 ( .A(data_valid), .Z(n148) );
  GTECH_AND2 U233 ( .A(n161), .B(n213), .Z(N222) );
  GTECH_NOT U234 ( .A(n204), .Z(n213) );
  GTECH_NOT U235 ( .A(n192), .Z(n161) );
  GTECH_NAND2 U236 ( .A(n211), .B(n177), .Z(n192) );
  GTECH_NOT U237 ( .A(n208), .Z(n211) );
  GTECH_OAI21 U238 ( .A(n196), .B(n203), .C(n214), .Z(N209) );
  GTECH_OR3 U239 ( .A(temp[17]), .B(n208), .C(n204), .Z(n214) );
  GTECH_NAND2 U240 ( .A(n215), .B(n216), .Z(n204) );
  GTECH_NOT U241 ( .A(n150), .Z(n215) );
  GTECH_NAND2 U242 ( .A(n162), .B(n157), .Z(n150) );
  GTECH_NOT U243 ( .A(n149), .Z(n162) );
  GTECH_NAND2 U244 ( .A(n206), .B(data_valid), .Z(n149) );
  GTECH_NAND2 U245 ( .A(data_valid), .B(n216), .Z(n203) );
  GTECH_NAND4 U246 ( .A(n217), .B(n199), .C(n153), .D(n182), .Z(n216) );
  GTECH_NAND2 U247 ( .A(n201), .B(n173), .Z(n182) );
  GTECH_NOT U248 ( .A(n218), .Z(n201) );
  GTECH_NAND2 U249 ( .A(temp[17]), .B(n177), .Z(n218) );
  GTECH_NAND4 U250 ( .A(temp[19]), .B(n206), .C(n187), .D(n157), .Z(n153) );
  GTECH_NOT U251 ( .A(temp[21]), .Z(n157) );
  GTECH_NOT U252 ( .A(n219), .Z(n206) );
  GTECH_OR3 U253 ( .A(n220), .B(n186), .C(n174), .Z(n199) );
  GTECH_NOT U254 ( .A(temp[16]), .Z(n174) );
  GTECH_NAND2 U255 ( .A(n180), .B(n177), .Z(n186) );
  GTECH_NOT U256 ( .A(temp[18]), .Z(n177) );
  GTECH_NOT U257 ( .A(temp[17]), .Z(n180) );
  GTECH_NOT U258 ( .A(n155), .Z(n217) );
  GTECH_OR3 U259 ( .A(temp[21]), .B(n221), .C(n219), .Z(n155) );
  GTECH_NAND2 U260 ( .A(n179), .B(n158), .Z(n219) );
  GTECH_NOT U261 ( .A(temp[22]), .Z(n179) );
  GTECH_NOT U262 ( .A(n196), .Z(n221) );
  GTECH_NAND2 U263 ( .A(temp[18]), .B(n173), .Z(n196) );
  GTECH_NOT U264 ( .A(n220), .Z(n173) );
  GTECH_NAND2 U265 ( .A(n222), .B(n158), .Z(n220) );
  GTECH_NOT U266 ( .A(temp[23]), .Z(n158) );
  GTECH_NOT U267 ( .A(n202), .Z(n222) );
  GTECH_OR3 U268 ( .A(temp[22]), .B(temp[21]), .C(n208), .Z(n202) );
  GTECH_NAND2 U269 ( .A(n223), .B(n187), .Z(n208) );
  GTECH_NOT U270 ( .A(temp[20]), .Z(n187) );
  GTECH_NOT U271 ( .A(temp[19]), .Z(n223) );
endmodule

