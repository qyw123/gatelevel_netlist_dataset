
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133;

  GTECH_XOR2 U86 ( .A(n67), .B(n68), .Z(sum[9]) );
  GTECH_XOR2 U87 ( .A(n69), .B(n70), .Z(sum[8]) );
  GTECH_XOR2 U88 ( .A(n71), .B(n72), .Z(sum[7]) );
  GTECH_OA21 U89 ( .A(n73), .B(n74), .C(n75), .Z(n72) );
  GTECH_XOR2 U90 ( .A(n74), .B(n73), .Z(sum[6]) );
  GTECH_OA21 U91 ( .A(n76), .B(n77), .C(n78), .Z(n73) );
  GTECH_XOR2 U92 ( .A(n77), .B(n76), .Z(sum[5]) );
  GTECH_OA21 U93 ( .A(n79), .B(n80), .C(n81), .Z(n76) );
  GTECH_XOR2 U94 ( .A(n80), .B(n79), .Z(sum[4]) );
  GTECH_XOR2 U95 ( .A(n82), .B(n83), .Z(sum[3]) );
  GTECH_OA21 U96 ( .A(n84), .B(n85), .C(n86), .Z(n83) );
  GTECH_XOR2 U97 ( .A(n85), .B(n84), .Z(sum[2]) );
  GTECH_OA21 U98 ( .A(n87), .B(n88), .C(n89), .Z(n84) );
  GTECH_XOR2 U99 ( .A(n88), .B(n87), .Z(sum[1]) );
  GTECH_OA21 U100 ( .A(n90), .B(n91), .C(n92), .Z(n87) );
  GTECH_XOR2 U101 ( .A(n93), .B(n94), .Z(sum[15]) );
  GTECH_AO21 U102 ( .A(n95), .B(n96), .C(n97), .Z(n93) );
  GTECH_XOR2 U103 ( .A(n95), .B(n96), .Z(sum[14]) );
  GTECH_AO21 U104 ( .A(n98), .B(n99), .C(n100), .Z(n95) );
  GTECH_XOR2 U105 ( .A(n99), .B(n98), .Z(sum[13]) );
  GTECH_AO21 U106 ( .A(cout), .B(n101), .C(n102), .Z(n98) );
  GTECH_XOR2 U107 ( .A(cout), .B(n101), .Z(sum[12]) );
  GTECH_XNOR2 U108 ( .A(n103), .B(n104), .Z(sum[11]) );
  GTECH_OAI21 U109 ( .A(n105), .B(n106), .C(n107), .Z(n103) );
  GTECH_XOR2 U110 ( .A(n106), .B(n105), .Z(sum[10]) );
  GTECH_OA21 U111 ( .A(n68), .B(n67), .C(n108), .Z(n105) );
  GTECH_OA21 U112 ( .A(n70), .B(n69), .C(n109), .Z(n68) );
  GTECH_XNOR2 U113 ( .A(cin), .B(n90), .Z(sum[0]) );
  GTECH_OAI21 U114 ( .A(n70), .B(n110), .C(n111), .Z(cout) );
  GTECH_OA21 U115 ( .A(n79), .B(n112), .C(n113), .Z(n70) );
  GTECH_OA21 U116 ( .A(n114), .B(n91), .C(n115), .Z(n79) );
  GTECH_NOT U117 ( .A(cin), .Z(n91) );
  GTECH_NOR3 U118 ( .A(n112), .B(n114), .C(n110), .Z(Pm) );
  GTECH_OR5 U119 ( .A(n88), .B(n82), .C(n85), .D(n90), .E(n116), .Z(n114) );
  GTECH_OAI21 U120 ( .A(b[0]), .B(a[0]), .C(n92), .Z(n90) );
  GTECH_OAI21 U121 ( .A(n117), .B(n110), .C(n111), .Z(Gm) );
  GTECH_AOI21 U122 ( .A(n118), .B(n94), .C(n119), .Z(n111) );
  GTECH_AO21 U123 ( .A(n120), .B(n96), .C(n97), .Z(n118) );
  GTECH_AO21 U124 ( .A(n99), .B(n102), .C(n100), .Z(n120) );
  GTECH_NAND4 U125 ( .A(n101), .B(n94), .C(n96), .D(n99), .Z(n110) );
  GTECH_OA21 U126 ( .A(b[13]), .B(a[13]), .C(n121), .Z(n99) );
  GTECH_NOT U127 ( .A(n100), .Z(n121) );
  GTECH_AND2 U128 ( .A(a[13]), .B(b[13]), .Z(n100) );
  GTECH_OA21 U129 ( .A(a[14]), .B(b[14]), .C(n122), .Z(n96) );
  GTECH_NOT U130 ( .A(n97), .Z(n122) );
  GTECH_AND2 U131 ( .A(a[14]), .B(b[14]), .Z(n97) );
  GTECH_OA21 U132 ( .A(a[15]), .B(b[15]), .C(n123), .Z(n94) );
  GTECH_NOT U133 ( .A(n119), .Z(n123) );
  GTECH_AND2 U134 ( .A(a[15]), .B(b[15]), .Z(n119) );
  GTECH_OA21 U135 ( .A(a[12]), .B(b[12]), .C(n124), .Z(n101) );
  GTECH_NOT U136 ( .A(n102), .Z(n124) );
  GTECH_AND2 U137 ( .A(a[12]), .B(b[12]), .Z(n102) );
  GTECH_OA21 U138 ( .A(n115), .B(n112), .C(n113), .Z(n117) );
  GTECH_OA21 U139 ( .A(n125), .B(n104), .C(n126), .Z(n113) );
  GTECH_OA21 U140 ( .A(n127), .B(n106), .C(n107), .Z(n125) );
  GTECH_OA21 U141 ( .A(n109), .B(n67), .C(n108), .Z(n127) );
  GTECH_OR4 U142 ( .A(n69), .B(n104), .C(n106), .D(n67), .Z(n112) );
  GTECH_OAI21 U143 ( .A(b[9]), .B(a[9]), .C(n108), .Z(n67) );
  GTECH_NAND2 U144 ( .A(a[9]), .B(b[9]), .Z(n108) );
  GTECH_OAI21 U145 ( .A(b[10]), .B(a[10]), .C(n107), .Z(n106) );
  GTECH_NAND2 U146 ( .A(b[10]), .B(a[10]), .Z(n107) );
  GTECH_OAI21 U147 ( .A(b[11]), .B(a[11]), .C(n126), .Z(n104) );
  GTECH_NAND2 U148 ( .A(a[11]), .B(b[11]), .Z(n126) );
  GTECH_OAI21 U149 ( .A(b[8]), .B(a[8]), .C(n109), .Z(n69) );
  GTECH_NAND2 U150 ( .A(a[8]), .B(b[8]), .Z(n109) );
  GTECH_AOI21 U151 ( .A(b[7]), .B(a[7]), .C(n128), .Z(n115) );
  GTECH_OAI22 U152 ( .A(n129), .B(n116), .C(n130), .D(n71), .Z(n128) );
  GTECH_OA21 U153 ( .A(n131), .B(n74), .C(n75), .Z(n130) );
  GTECH_OA21 U154 ( .A(n77), .B(n81), .C(n78), .Z(n131) );
  GTECH_OR4 U155 ( .A(n80), .B(n74), .C(n77), .D(n71), .Z(n116) );
  GTECH_XNOR2 U156 ( .A(a[7]), .B(b[7]), .Z(n71) );
  GTECH_OAI21 U157 ( .A(b[5]), .B(a[5]), .C(n78), .Z(n77) );
  GTECH_NAND2 U158 ( .A(b[5]), .B(a[5]), .Z(n78) );
  GTECH_OAI21 U159 ( .A(b[6]), .B(a[6]), .C(n75), .Z(n74) );
  GTECH_NAND2 U160 ( .A(b[6]), .B(a[6]), .Z(n75) );
  GTECH_OAI21 U161 ( .A(b[4]), .B(a[4]), .C(n81), .Z(n80) );
  GTECH_NAND2 U162 ( .A(b[4]), .B(a[4]), .Z(n81) );
  GTECH_AOI2N2 U163 ( .A(b[3]), .B(a[3]), .C(n132), .D(n82), .Z(n129) );
  GTECH_XNOR2 U164 ( .A(a[3]), .B(b[3]), .Z(n82) );
  GTECH_OA21 U165 ( .A(n133), .B(n85), .C(n86), .Z(n132) );
  GTECH_OAI21 U166 ( .A(b[2]), .B(a[2]), .C(n86), .Z(n85) );
  GTECH_NAND2 U167 ( .A(b[2]), .B(a[2]), .Z(n86) );
  GTECH_OA21 U168 ( .A(n92), .B(n88), .C(n89), .Z(n133) );
  GTECH_OAI21 U169 ( .A(b[1]), .B(a[1]), .C(n89), .Z(n88) );
  GTECH_NAND2 U170 ( .A(b[1]), .B(a[1]), .Z(n89) );
  GTECH_NAND2 U171 ( .A(a[0]), .B(b[0]), .Z(n92) );
endmodule

