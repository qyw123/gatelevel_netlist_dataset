
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384;

  GTECH_OAI22 U140 ( .A(n279), .B(n280), .C(n281), .D(n282), .Z(sum[9]) );
  GTECH_XOR2 U141 ( .A(n283), .B(n284), .Z(n281) );
  GTECH_XOR2 U142 ( .A(n285), .B(n283), .Z(n280) );
  GTECH_OAI21 U143 ( .A(a[9]), .B(b[9]), .C(n286), .Z(n283) );
  GTECH_NOT U144 ( .A(n287), .Z(n286) );
  GTECH_AO21 U145 ( .A(n288), .B(n279), .C(n289), .Z(sum[8]) );
  GTECH_OAI22 U146 ( .A(n290), .B(n291), .C(n292), .D(n293), .Z(sum[7]) );
  GTECH_XNOR2 U147 ( .A(n294), .B(n295), .Z(n292) );
  GTECH_XOR2 U148 ( .A(n296), .B(n295), .Z(n290) );
  GTECH_XOR2 U149 ( .A(a[7]), .B(b[7]), .Z(n295) );
  GTECH_OA21 U150 ( .A(n297), .B(n298), .C(n299), .Z(n296) );
  GTECH_OAI22 U151 ( .A(n300), .B(n291), .C(n301), .D(n293), .Z(sum[6]) );
  GTECH_XNOR2 U152 ( .A(n302), .B(n303), .Z(n301) );
  GTECH_XNOR2 U153 ( .A(n303), .B(n298), .Z(n300) );
  GTECH_AOI21 U154 ( .A(n304), .B(n305), .C(n306), .Z(n298) );
  GTECH_OR_NOT U155 ( .A(n297), .B(n299), .Z(n303) );
  GTECH_OAI2N2 U156 ( .A(n307), .B(n308), .C(n309), .D(n307), .Z(sum[5]) );
  GTECH_OAI21 U157 ( .A(n305), .B(n291), .C(n310), .Z(n309) );
  GTECH_AOI21 U158 ( .A(n310), .B(n291), .C(n305), .Z(n308) );
  GTECH_AND2 U159 ( .A(n311), .B(n304), .Z(n307) );
  GTECH_NOT U160 ( .A(n306), .Z(n311) );
  GTECH_XNOR2 U161 ( .A(n291), .B(n312), .Z(sum[4]) );
  GTECH_OAI22 U162 ( .A(n313), .B(n314), .C(cin), .D(n315), .Z(sum[3]) );
  GTECH_XOR2 U163 ( .A(n316), .B(n317), .Z(n315) );
  GTECH_OA21 U164 ( .A(n318), .B(n319), .C(n320), .Z(n316) );
  GTECH_XNOR2 U165 ( .A(n321), .B(n317), .Z(n314) );
  GTECH_XOR2 U166 ( .A(a[3]), .B(b[3]), .Z(n317) );
  GTECH_OAI22 U167 ( .A(n313), .B(n322), .C(cin), .D(n323), .Z(sum[2]) );
  GTECH_XNOR2 U168 ( .A(n324), .B(n319), .Z(n323) );
  GTECH_AOI21 U169 ( .A(n325), .B(n326), .C(n327), .Z(n319) );
  GTECH_XNOR2 U170 ( .A(n328), .B(n324), .Z(n322) );
  GTECH_OR_NOT U171 ( .A(n318), .B(n320), .Z(n324) );
  GTECH_OAI2N2 U172 ( .A(n329), .B(n330), .C(n331), .D(n329), .Z(sum[1]) );
  GTECH_OAI21 U173 ( .A(cin), .B(n326), .C(n332), .Z(n331) );
  GTECH_AOI21 U174 ( .A(n332), .B(cin), .C(n326), .Z(n330) );
  GTECH_AND2 U175 ( .A(a[0]), .B(b[0]), .Z(n326) );
  GTECH_AND2 U176 ( .A(n333), .B(n325), .Z(n329) );
  GTECH_NOT U177 ( .A(n327), .Z(n333) );
  GTECH_OAI22 U178 ( .A(n334), .B(n335), .C(n336), .D(n337), .Z(sum[15]) );
  GTECH_XNOR2 U179 ( .A(n338), .B(n339), .Z(n337) );
  GTECH_XOR2 U180 ( .A(n340), .B(n339), .Z(n335) );
  GTECH_XOR2 U181 ( .A(a[15]), .B(b[15]), .Z(n339) );
  GTECH_OA21 U182 ( .A(n341), .B(n342), .C(n343), .Z(n340) );
  GTECH_OAI22 U183 ( .A(n334), .B(n344), .C(n336), .D(n345), .Z(sum[14]) );
  GTECH_XNOR2 U184 ( .A(n346), .B(n347), .Z(n345) );
  GTECH_XNOR2 U185 ( .A(n347), .B(n341), .Z(n344) );
  GTECH_AOI21 U186 ( .A(n348), .B(n349), .C(n350), .Z(n341) );
  GTECH_NOT U187 ( .A(n351), .Z(n348) );
  GTECH_OR_NOT U188 ( .A(n342), .B(n343), .Z(n347) );
  GTECH_OAI22 U189 ( .A(n334), .B(n352), .C(n336), .D(n353), .Z(sum[13]) );
  GTECH_XNOR2 U190 ( .A(n354), .B(n355), .Z(n353) );
  GTECH_XOR2 U191 ( .A(n355), .B(n356), .Z(n352) );
  GTECH_NOR2 U192 ( .A(n350), .B(n351), .Z(n355) );
  GTECH_NAND2 U193 ( .A(n357), .B(n358), .Z(sum[12]) );
  GTECH_OAI21 U194 ( .A(n349), .B(n359), .C(n334), .Z(n358) );
  GTECH_NOT U195 ( .A(n336), .Z(n334) );
  GTECH_OAI22 U196 ( .A(n360), .B(n279), .C(n361), .D(n282), .Z(sum[11]) );
  GTECH_XNOR2 U197 ( .A(n362), .B(n363), .Z(n361) );
  GTECH_XOR2 U198 ( .A(n364), .B(n363), .Z(n360) );
  GTECH_XOR2 U199 ( .A(a[11]), .B(b[11]), .Z(n363) );
  GTECH_OA21 U200 ( .A(n365), .B(n366), .C(n367), .Z(n364) );
  GTECH_NOT U201 ( .A(n368), .Z(n367) );
  GTECH_OAI22 U202 ( .A(n282), .B(n369), .C(n279), .D(n370), .Z(sum[10]) );
  GTECH_XOR2 U203 ( .A(n366), .B(n371), .Z(n370) );
  GTECH_OAI21 U204 ( .A(n287), .B(n285), .C(n372), .Z(n366) );
  GTECH_XNOR2 U205 ( .A(n373), .B(n371), .Z(n369) );
  GTECH_NOR2 U206 ( .A(n365), .B(n368), .Z(n371) );
  GTECH_NOT U207 ( .A(n279), .Z(n282) );
  GTECH_XNOR2 U208 ( .A(n313), .B(n374), .Z(sum[0]) );
  GTECH_OAI21 U209 ( .A(n336), .B(n375), .C(n357), .Z(cout) );
  GTECH_NAND3 U210 ( .A(n354), .B(n356), .C(n336), .Z(n357) );
  GTECH_NOT U211 ( .A(n349), .Z(n356) );
  GTECH_AND2 U212 ( .A(b[12]), .B(a[12]), .Z(n349) );
  GTECH_AOI21 U213 ( .A(n338), .B(a[15]), .C(n376), .Z(n375) );
  GTECH_OA21 U214 ( .A(a[15]), .B(n338), .C(b[15]), .Z(n376) );
  GTECH_OAI21 U215 ( .A(n346), .B(n342), .C(n343), .Z(n338) );
  GTECH_NAND2 U216 ( .A(a[14]), .B(b[14]), .Z(n343) );
  GTECH_NOR2 U217 ( .A(b[14]), .B(a[14]), .Z(n342) );
  GTECH_OA21 U218 ( .A(n351), .B(n359), .C(n377), .Z(n346) );
  GTECH_NOT U219 ( .A(n350), .Z(n377) );
  GTECH_AND2 U220 ( .A(a[13]), .B(b[13]), .Z(n350) );
  GTECH_NOT U221 ( .A(n354), .Z(n359) );
  GTECH_OR2 U222 ( .A(b[12]), .B(a[12]), .Z(n354) );
  GTECH_NOR2 U223 ( .A(a[13]), .B(b[13]), .Z(n351) );
  GTECH_AOI21 U224 ( .A(n279), .B(n378), .C(n289), .Z(n336) );
  GTECH_NOR2 U225 ( .A(n288), .B(n279), .Z(n289) );
  GTECH_OR_NOT U226 ( .A(n285), .B(n284), .Z(n288) );
  GTECH_AND2 U227 ( .A(b[8]), .B(a[8]), .Z(n285) );
  GTECH_OA21 U228 ( .A(a[11]), .B(n362), .C(n379), .Z(n378) );
  GTECH_AO21 U229 ( .A(n362), .B(a[11]), .C(b[11]), .Z(n379) );
  GTECH_AO21 U230 ( .A(n380), .B(n373), .C(n368), .Z(n362) );
  GTECH_AND2 U231 ( .A(b[10]), .B(a[10]), .Z(n368) );
  GTECH_OA21 U232 ( .A(n287), .B(n284), .C(n372), .Z(n373) );
  GTECH_OR2 U233 ( .A(a[9]), .B(b[9]), .Z(n372) );
  GTECH_OR2 U234 ( .A(b[8]), .B(a[8]), .Z(n284) );
  GTECH_AND2 U235 ( .A(b[9]), .B(a[9]), .Z(n287) );
  GTECH_NOT U236 ( .A(n365), .Z(n380) );
  GTECH_NOR2 U237 ( .A(b[10]), .B(a[10]), .Z(n365) );
  GTECH_OAI22 U238 ( .A(n291), .B(n312), .C(n381), .D(n293), .Z(n279) );
  GTECH_AOI21 U239 ( .A(n294), .B(a[7]), .C(n382), .Z(n381) );
  GTECH_OA21 U240 ( .A(a[7]), .B(n294), .C(b[7]), .Z(n382) );
  GTECH_OAI21 U241 ( .A(n302), .B(n297), .C(n299), .Z(n294) );
  GTECH_NAND2 U242 ( .A(a[6]), .B(b[6]), .Z(n299) );
  GTECH_NOR2 U243 ( .A(b[6]), .B(a[6]), .Z(n297) );
  GTECH_AOI21 U244 ( .A(n304), .B(n310), .C(n306), .Z(n302) );
  GTECH_AND2 U245 ( .A(a[5]), .B(b[5]), .Z(n306) );
  GTECH_OR2 U246 ( .A(a[5]), .B(b[5]), .Z(n304) );
  GTECH_OR_NOT U247 ( .A(n305), .B(n310), .Z(n312) );
  GTECH_OR2 U248 ( .A(a[4]), .B(b[4]), .Z(n310) );
  GTECH_AND2 U249 ( .A(b[4]), .B(a[4]), .Z(n305) );
  GTECH_NOT U250 ( .A(n293), .Z(n291) );
  GTECH_AOI2N2 U251 ( .A(n313), .B(n374), .C(n383), .D(n313), .Z(n293) );
  GTECH_AOI21 U252 ( .A(n321), .B(a[3]), .C(n384), .Z(n383) );
  GTECH_OA21 U253 ( .A(a[3]), .B(n321), .C(b[3]), .Z(n384) );
  GTECH_OAI21 U254 ( .A(n328), .B(n318), .C(n320), .Z(n321) );
  GTECH_NAND2 U255 ( .A(a[2]), .B(b[2]), .Z(n320) );
  GTECH_NOR2 U256 ( .A(b[2]), .B(a[2]), .Z(n318) );
  GTECH_AOI21 U257 ( .A(n325), .B(n332), .C(n327), .Z(n328) );
  GTECH_AND2 U258 ( .A(a[1]), .B(b[1]), .Z(n327) );
  GTECH_OR2 U259 ( .A(b[0]), .B(a[0]), .Z(n332) );
  GTECH_OR2 U260 ( .A(a[1]), .B(b[1]), .Z(n325) );
  GTECH_XOR2 U261 ( .A(a[0]), .B(b[0]), .Z(n374) );
  GTECH_NOT U262 ( .A(cin), .Z(n313) );
endmodule

