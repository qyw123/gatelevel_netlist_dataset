
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131;

  GTECH_XOR2 U86 ( .A(n67), .B(n68), .Z(sum[9]) );
  GTECH_XOR2 U87 ( .A(n69), .B(n70), .Z(sum[8]) );
  GTECH_XNOR2 U88 ( .A(n71), .B(n72), .Z(sum[7]) );
  GTECH_AOI21 U89 ( .A(n73), .B(n74), .C(n75), .Z(n72) );
  GTECH_XOR2 U90 ( .A(n74), .B(n73), .Z(sum[6]) );
  GTECH_AO22 U91 ( .A(b[5]), .B(a[5]), .C(n76), .D(n77), .Z(n73) );
  GTECH_XOR2 U92 ( .A(n77), .B(n76), .Z(sum[5]) );
  GTECH_AO22 U93 ( .A(b[4]), .B(a[4]), .C(n78), .D(n79), .Z(n76) );
  GTECH_XOR2 U94 ( .A(n79), .B(n78), .Z(sum[4]) );
  GTECH_NOT U95 ( .A(n80), .Z(n78) );
  GTECH_XNOR2 U96 ( .A(n81), .B(n82), .Z(sum[3]) );
  GTECH_AOI21 U97 ( .A(n83), .B(n84), .C(n85), .Z(n82) );
  GTECH_XOR2 U98 ( .A(n84), .B(n83), .Z(sum[2]) );
  GTECH_AO22 U99 ( .A(b[1]), .B(a[1]), .C(n86), .D(n87), .Z(n83) );
  GTECH_XOR2 U100 ( .A(n87), .B(n86), .Z(sum[1]) );
  GTECH_AO22 U101 ( .A(a[0]), .B(b[0]), .C(n88), .D(cin), .Z(n86) );
  GTECH_XNOR2 U102 ( .A(n89), .B(n90), .Z(sum[15]) );
  GTECH_AOI21 U103 ( .A(n91), .B(n92), .C(n93), .Z(n90) );
  GTECH_XOR2 U104 ( .A(n92), .B(n91), .Z(sum[14]) );
  GTECH_AO21 U105 ( .A(n94), .B(n95), .C(n96), .Z(n91) );
  GTECH_XOR2 U106 ( .A(n94), .B(n95), .Z(sum[13]) );
  GTECH_AO22 U107 ( .A(a[12]), .B(b[12]), .C(cout), .D(n97), .Z(n94) );
  GTECH_XOR2 U108 ( .A(n97), .B(cout), .Z(sum[12]) );
  GTECH_XOR2 U109 ( .A(n98), .B(n99), .Z(sum[11]) );
  GTECH_OA21 U110 ( .A(n100), .B(n101), .C(n102), .Z(n99) );
  GTECH_XOR2 U111 ( .A(n101), .B(n100), .Z(sum[10]) );
  GTECH_OA21 U112 ( .A(n67), .B(n68), .C(n103), .Z(n100) );
  GTECH_OA21 U113 ( .A(n70), .B(n69), .C(n104), .Z(n67) );
  GTECH_XNOR2 U114 ( .A(n105), .B(n88), .Z(sum[0]) );
  GTECH_OAI21 U115 ( .A(n70), .B(n106), .C(n107), .Z(cout) );
  GTECH_OA21 U116 ( .A(n80), .B(n108), .C(n109), .Z(n70) );
  GTECH_OA21 U117 ( .A(n110), .B(n105), .C(n111), .Z(n80) );
  GTECH_NOT U118 ( .A(cin), .Z(n105) );
  GTECH_NOR3 U119 ( .A(n108), .B(n110), .C(n106), .Z(Pm) );
  GTECH_NAND5 U120 ( .A(n84), .B(n87), .C(n81), .D(n112), .E(n88), .Z(n110) );
  GTECH_XOR2 U121 ( .A(a[0]), .B(b[0]), .Z(n88) );
  GTECH_OAI21 U122 ( .A(n113), .B(n106), .C(n107), .Z(Gm) );
  GTECH_AOI21 U123 ( .A(b[15]), .B(a[15]), .C(n114), .Z(n107) );
  GTECH_OA21 U124 ( .A(n93), .B(n115), .C(n89), .Z(n114) );
  GTECH_OA21 U125 ( .A(n116), .B(n96), .C(n92), .Z(n115) );
  GTECH_NOT U126 ( .A(n117), .Z(n96) );
  GTECH_AND3 U127 ( .A(a[12]), .B(n95), .C(b[12]), .Z(n116) );
  GTECH_NOT U128 ( .A(n118), .Z(n93) );
  GTECH_NAND4 U129 ( .A(n92), .B(n95), .C(n97), .D(n89), .Z(n106) );
  GTECH_XOR2 U130 ( .A(a[15]), .B(b[15]), .Z(n89) );
  GTECH_XOR2 U131 ( .A(a[12]), .B(b[12]), .Z(n97) );
  GTECH_OA21 U132 ( .A(b[13]), .B(a[13]), .C(n117), .Z(n95) );
  GTECH_NAND2 U133 ( .A(a[13]), .B(b[13]), .Z(n117) );
  GTECH_OA21 U134 ( .A(b[14]), .B(a[14]), .C(n118), .Z(n92) );
  GTECH_NAND2 U135 ( .A(a[14]), .B(b[14]), .Z(n118) );
  GTECH_OA21 U136 ( .A(n111), .B(n108), .C(n109), .Z(n113) );
  GTECH_AOI2N2 U137 ( .A(b[11]), .B(a[11]), .C(n119), .D(n98), .Z(n109) );
  GTECH_OA21 U138 ( .A(n120), .B(n101), .C(n102), .Z(n119) );
  GTECH_NAND2 U139 ( .A(a[10]), .B(b[10]), .Z(n102) );
  GTECH_OA21 U140 ( .A(n104), .B(n68), .C(n103), .Z(n120) );
  GTECH_NAND2 U141 ( .A(b[8]), .B(a[8]), .Z(n104) );
  GTECH_OR4 U142 ( .A(n68), .B(n69), .C(n98), .D(n101), .Z(n108) );
  GTECH_XNOR2 U143 ( .A(a[10]), .B(b[10]), .Z(n101) );
  GTECH_XNOR2 U144 ( .A(a[11]), .B(b[11]), .Z(n98) );
  GTECH_XNOR2 U145 ( .A(a[8]), .B(b[8]), .Z(n69) );
  GTECH_OAI21 U146 ( .A(a[9]), .B(b[9]), .C(n103), .Z(n68) );
  GTECH_NAND2 U147 ( .A(b[9]), .B(a[9]), .Z(n103) );
  GTECH_AOI222 U148 ( .A(a[7]), .B(b[7]), .C(n112), .D(n121), .E(n71), .F(n122), .Z(n111) );
  GTECH_AO21 U149 ( .A(n123), .B(n74), .C(n75), .Z(n122) );
  GTECH_AND2 U150 ( .A(a[6]), .B(b[6]), .Z(n75) );
  GTECH_AO21 U151 ( .A(b[5]), .B(a[5]), .C(n124), .Z(n123) );
  GTECH_NOT U152 ( .A(n125), .Z(n124) );
  GTECH_NAND3 U153 ( .A(b[4]), .B(n77), .C(a[4]), .Z(n125) );
  GTECH_AO22 U154 ( .A(b[3]), .B(a[3]), .C(n126), .D(n81), .Z(n121) );
  GTECH_XOR2 U155 ( .A(a[3]), .B(b[3]), .Z(n81) );
  GTECH_AO21 U156 ( .A(n127), .B(n84), .C(n85), .Z(n126) );
  GTECH_AND2 U157 ( .A(a[2]), .B(b[2]), .Z(n85) );
  GTECH_XOR2 U158 ( .A(a[2]), .B(b[2]), .Z(n84) );
  GTECH_AO21 U159 ( .A(b[1]), .B(a[1]), .C(n128), .Z(n127) );
  GTECH_NOT U160 ( .A(n129), .Z(n128) );
  GTECH_NAND3 U161 ( .A(a[0]), .B(n87), .C(b[0]), .Z(n129) );
  GTECH_XNOR2 U162 ( .A(a[1]), .B(n130), .Z(n87) );
  GTECH_NOT U163 ( .A(b[1]), .Z(n130) );
  GTECH_AND4 U164 ( .A(n79), .B(n77), .C(n74), .D(n71), .Z(n112) );
  GTECH_XOR2 U165 ( .A(a[7]), .B(b[7]), .Z(n71) );
  GTECH_XOR2 U166 ( .A(a[6]), .B(b[6]), .Z(n74) );
  GTECH_XNOR2 U167 ( .A(a[5]), .B(n131), .Z(n77) );
  GTECH_NOT U168 ( .A(b[5]), .Z(n131) );
  GTECH_XOR2 U169 ( .A(a[4]), .B(b[4]), .Z(n79) );
endmodule

