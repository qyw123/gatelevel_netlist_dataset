
module CRC_16_parallel ( clk, rst_n, data, data_valid, crc );
  input [7:0] data;
  output [15:0] crc;
  input clk, rst_n, data_valid;
  wire   N11, N15, N23, N34, N37, N39, N41, N43, N45, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N58, N60, N62, N64, N69, N70, N99, N209,
         N222, N235, N248, N261, N274, N287, N298, N307, N316, N323, N328,
         N331, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229;
  wire   [23:0] temp;

  GTECH_FJK2S temp_reg_15_ ( .J(n106), .K(n106), .TI(N56), .TE(N287), .CP(clk), 
        .CD(rst_n), .Q(temp[15]) );
  GTECH_FJK2S temp_reg_14_ ( .J(n106), .K(n106), .TI(N55), .TE(N209), .CP(clk), 
        .CD(rst_n), .Q(temp[14]) );
  GTECH_FJK2S temp_reg_13_ ( .J(n106), .K(n106), .TI(N54), .TE(N222), .CP(clk), 
        .CD(rst_n), .Q(temp[13]) );
  GTECH_FJK2S temp_reg_12_ ( .J(n106), .K(n106), .TI(N53), .TE(N235), .CP(clk), 
        .CD(rst_n), .Q(temp[12]), .QN(N53) );
  GTECH_FJK2S temp_reg_11_ ( .J(n106), .K(n106), .TI(N52), .TE(N248), .CP(clk), 
        .CD(rst_n), .Q(temp[11]) );
  GTECH_FJK2S temp_reg_10_ ( .J(n106), .K(n106), .TI(N51), .TE(N261), .CP(clk), 
        .CD(rst_n), .Q(temp[10]) );
  GTECH_FJK2S temp_reg_9_ ( .J(n106), .K(n106), .TI(N50), .TE(N274), .CP(clk), 
        .CD(rst_n), .Q(temp[9]) );
  GTECH_FJK2S temp_reg_8_ ( .J(n106), .K(n106), .TI(N49), .TE(N287), .CP(clk), 
        .CD(rst_n), .Q(temp[8]) );
  GTECH_FJK2S temp_reg_7_ ( .J(n106), .K(n106), .TI(N48), .TE(N298), .CP(clk), 
        .CD(rst_n), .Q(temp[7]) );
  GTECH_FJK2S temp_reg_6_ ( .J(n106), .K(n106), .TI(N47), .TE(N307), .CP(clk), 
        .CD(rst_n), .Q(temp[6]) );
  GTECH_FJK2S temp_reg_5_ ( .J(n106), .K(n106), .TI(N45), .TE(N316), .CP(clk), 
        .CD(rst_n), .Q(temp[5]), .QN(N45) );
  GTECH_FJK2S temp_reg_4_ ( .J(n106), .K(n106), .TI(N43), .TE(N323), .CP(clk), 
        .CD(rst_n), .Q(temp[4]) );
  GTECH_FJK2S temp_reg_3_ ( .J(n106), .K(n106), .TI(N41), .TE(N328), .CP(clk), 
        .CD(rst_n), .Q(temp[3]) );
  GTECH_FJK2S temp_reg_2_ ( .J(n106), .K(n106), .TI(N39), .TE(N331), .CP(clk), 
        .CD(rst_n), .Q(temp[2]) );
  GTECH_FJK2S temp_reg_1_ ( .J(n106), .K(n106), .TI(N37), .TE(N70), .CP(clk), 
        .CD(rst_n), .Q(temp[1]) );
  GTECH_FJK2S temp_reg_0_ ( .J(n106), .K(n106), .TI(N34), .TE(N69), .CP(clk), 
        .CD(rst_n), .Q(temp[0]), .QN(N34) );
  GTECH_FJK2S crc_reg_15_ ( .J(n106), .K(n106), .TI(temp[15]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[15]) );
  GTECH_FJK2S crc_reg_14_ ( .J(n106), .K(n106), .TI(temp[14]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[14]) );
  GTECH_FJK2S crc_reg_13_ ( .J(n106), .K(n106), .TI(temp[13]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[13]) );
  GTECH_FJK2S crc_reg_12_ ( .J(n106), .K(n106), .TI(temp[12]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[12]) );
  GTECH_FJK2S crc_reg_11_ ( .J(n106), .K(n106), .TI(temp[11]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[11]) );
  GTECH_FJK2S crc_reg_10_ ( .J(n106), .K(n106), .TI(temp[10]), .TE(N99), .CP(
        clk), .CD(rst_n), .Q(crc[10]) );
  GTECH_FJK2S crc_reg_9_ ( .J(n106), .K(n106), .TI(temp[9]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[9]) );
  GTECH_FJK2S crc_reg_8_ ( .J(n106), .K(n106), .TI(temp[8]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[8]) );
  GTECH_FJK2S crc_reg_7_ ( .J(n106), .K(n106), .TI(temp[7]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[7]) );
  GTECH_FJK2S crc_reg_6_ ( .J(n106), .K(n106), .TI(temp[6]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[6]) );
  GTECH_FJK2S crc_reg_5_ ( .J(n106), .K(n106), .TI(temp[5]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[5]) );
  GTECH_FJK2S crc_reg_4_ ( .J(n106), .K(n106), .TI(temp[4]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[4]) );
  GTECH_FJK2S crc_reg_3_ ( .J(n106), .K(n106), .TI(temp[3]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[3]) );
  GTECH_FJK2S crc_reg_2_ ( .J(n106), .K(n106), .TI(temp[2]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[2]) );
  GTECH_FJK2S crc_reg_1_ ( .J(n106), .K(n106), .TI(temp[1]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[1]) );
  GTECH_FJK2S crc_reg_0_ ( .J(n106), .K(n106), .TI(temp[0]), .TE(N99), .CP(clk), .CD(rst_n), .Q(crc[0]) );
  GTECH_FD3 temp_reg_23_ ( .D(n105), .CP(clk), .CD(n97), .SD(n96), .Q(temp[23]), .QN(N11) );
  GTECH_FD3 temp_reg_22_ ( .D(n104), .CP(clk), .CD(n95), .SD(n94), .Q(temp[22]), .QN(N15) );
  GTECH_FD3 temp_reg_21_ ( .D(n103), .CP(clk), .CD(n93), .SD(n92), .Q(temp[21]) );
  GTECH_FD3 temp_reg_20_ ( .D(n102), .CP(clk), .CD(n91), .SD(n90), .Q(temp[20]), .QN(N23) );
  GTECH_FD3 temp_reg_19_ ( .D(n101), .CP(clk), .CD(n89), .SD(n88), .Q(temp[19]), .QN(N64) );
  GTECH_FD3 temp_reg_18_ ( .D(n100), .CP(clk), .CD(n87), .SD(n86), .Q(temp[18]), .QN(N62) );
  GTECH_FD3 temp_reg_17_ ( .D(n99), .CP(clk), .CD(n85), .SD(n84), .Q(temp[17]), 
        .QN(N60) );
  GTECH_FD3 temp_reg_16_ ( .D(n98), .CP(clk), .CD(n83), .SD(n82), .Q(temp[16]), 
        .QN(N58) );
  GTECH_ZERO U149 ( .Z(n106) );
  GTECH_MUX2 U150 ( .A(n154), .B(n155), .S(temp[17]), .Z(n99) );
  GTECH_OAI21 U151 ( .A(temp[21]), .B(n156), .C(n157), .Z(n155) );
  GTECH_AND2 U152 ( .A(temp[21]), .B(n157), .Z(n154) );
  GTECH_XOR2 U153 ( .A(N274), .B(temp[16]), .Z(n98) );
  GTECH_NAND2 U154 ( .A(n158), .B(n159), .Z(n97) );
  GTECH_NOT U155 ( .A(data[7]), .Z(n159) );
  GTECH_NAND2 U156 ( .A(data[7]), .B(n158), .Z(n96) );
  GTECH_NAND2 U157 ( .A(n158), .B(n160), .Z(n95) );
  GTECH_NOT U158 ( .A(data[6]), .Z(n160) );
  GTECH_NAND2 U159 ( .A(data[6]), .B(n158), .Z(n94) );
  GTECH_NAND2 U160 ( .A(n158), .B(n161), .Z(n93) );
  GTECH_NOT U161 ( .A(data[5]), .Z(n161) );
  GTECH_NAND2 U162 ( .A(data[5]), .B(n158), .Z(n92) );
  GTECH_NAND2 U163 ( .A(n158), .B(n162), .Z(n91) );
  GTECH_NOT U164 ( .A(data[4]), .Z(n162) );
  GTECH_NAND2 U165 ( .A(data[4]), .B(n158), .Z(n90) );
  GTECH_NAND2 U166 ( .A(n158), .B(n163), .Z(n89) );
  GTECH_NOT U167 ( .A(data[3]), .Z(n163) );
  GTECH_NAND2 U168 ( .A(data[3]), .B(n158), .Z(n88) );
  GTECH_NAND2 U169 ( .A(n158), .B(n164), .Z(n87) );
  GTECH_NOT U170 ( .A(data[2]), .Z(n164) );
  GTECH_NAND2 U171 ( .A(data[2]), .B(n158), .Z(n86) );
  GTECH_NAND2 U172 ( .A(n158), .B(n165), .Z(n85) );
  GTECH_NOT U173 ( .A(data[1]), .Z(n165) );
  GTECH_NAND2 U174 ( .A(data[1]), .B(n158), .Z(n84) );
  GTECH_NAND2 U175 ( .A(n158), .B(n166), .Z(n83) );
  GTECH_NOT U176 ( .A(data[0]), .Z(n166) );
  GTECH_NAND2 U177 ( .A(data[0]), .B(n158), .Z(n82) );
  GTECH_NOT U178 ( .A(rst_n), .Z(n158) );
  GTECH_AND2 U179 ( .A(temp[23]), .B(n167), .Z(n105) );
  GTECH_AOI21 U180 ( .A(data_valid), .B(n168), .C(n169), .Z(n104) );
  GTECH_AND2 U181 ( .A(temp[21]), .B(n170), .Z(n103) );
  GTECH_AND2 U182 ( .A(temp[20]), .B(n171), .Z(n102) );
  GTECH_XOR2 U183 ( .A(temp[19]), .B(n172), .Z(n101) );
  GTECH_AND3 U184 ( .A(n173), .B(n174), .C(data_valid), .Z(n172) );
  GTECH_NAND2 U185 ( .A(n175), .B(n176), .Z(n174) );
  GTECH_XOR2 U186 ( .A(temp[18]), .B(n177), .Z(n100) );
  GTECH_AND4 U187 ( .A(data_valid), .B(n178), .C(n179), .D(n168), .Z(n177) );
  GTECH_OAI21 U188 ( .A(temp[21]), .B(n180), .C(n169), .Z(n178) );
  GTECH_AND4 U189 ( .A(n181), .B(n182), .C(data_valid), .D(n183), .Z(N99) );
  GTECH_NOT U190 ( .A(temp[16]), .Z(n183) );
  GTECH_NOT U191 ( .A(n184), .Z(N69) );
  GTECH_XOR2 U192 ( .A(temp[19]), .B(temp[15]), .Z(N56) );
  GTECH_XOR2 U193 ( .A(temp[18]), .B(temp[14]), .Z(N55) );
  GTECH_XOR2 U194 ( .A(temp[17]), .B(temp[13]), .Z(N54) );
  GTECH_XOR2 U195 ( .A(temp[22]), .B(temp[11]), .Z(N52) );
  GTECH_XOR2 U196 ( .A(temp[21]), .B(temp[10]), .Z(N51) );
  GTECH_XOR2 U197 ( .A(temp[9]), .B(temp[20]), .Z(N50) );
  GTECH_XOR2 U198 ( .A(temp[8]), .B(temp[19]), .Z(N49) );
  GTECH_XOR2 U199 ( .A(n185), .B(temp[7]), .Z(N48) );
  GTECH_NAND2 U200 ( .A(n168), .B(n186), .Z(n185) );
  GTECH_XOR2 U201 ( .A(n187), .B(temp[6]), .Z(N47) );
  GTECH_NAND2 U202 ( .A(n169), .B(n188), .Z(n187) );
  GTECH_XOR2 U203 ( .A(temp[4]), .B(temp[20]), .Z(N43) );
  GTECH_XOR2 U204 ( .A(temp[3]), .B(temp[19]), .Z(N41) );
  GTECH_XOR2 U205 ( .A(temp[2]), .B(temp[18]), .Z(N39) );
  GTECH_XOR2 U206 ( .A(temp[1]), .B(temp[17]), .Z(N37) );
  GTECH_AND2 U207 ( .A(n189), .B(n190), .Z(N331) );
  GTECH_AOI21 U208 ( .A(n191), .B(n192), .C(n193), .Z(N328) );
  GTECH_AND2 U209 ( .A(n194), .B(n195), .Z(N323) );
  GTECH_OAI21 U210 ( .A(temp[19]), .B(n192), .C(n196), .Z(n194) );
  GTECH_AND2 U211 ( .A(n197), .B(n198), .Z(N316) );
  GTECH_OAI21 U212 ( .A(n170), .B(n199), .C(n200), .Z(n197) );
  GTECH_AND2 U213 ( .A(n201), .B(n202), .Z(N307) );
  GTECH_OAI21 U214 ( .A(n167), .B(n173), .C(n200), .Z(n202) );
  GTECH_NOT U215 ( .A(n195), .Z(n200) );
  GTECH_OAI21 U216 ( .A(n171), .B(n196), .C(n193), .Z(n195) );
  GTECH_AND_NOT U217 ( .A(n203), .B(n189), .Z(n193) );
  GTECH_OAI21 U218 ( .A(n167), .B(n204), .C(n205), .Z(n189) );
  GTECH_NOT U219 ( .A(N70), .Z(n205) );
  GTECH_OAI21 U220 ( .A(n167), .B(n190), .C(n184), .Z(N70) );
  GTECH_NAND2 U221 ( .A(n206), .B(data_valid), .Z(n184) );
  GTECH_NOT U222 ( .A(n207), .Z(n206) );
  GTECH_NAND3 U223 ( .A(data_valid), .B(n208), .C(n175), .Z(n203) );
  GTECH_NAND2 U224 ( .A(n168), .B(n209), .Z(n173) );
  GTECH_OAI21 U225 ( .A(temp[21]), .B(n210), .C(n157), .Z(n201) );
  GTECH_OAI22 U226 ( .A(n167), .B(n168), .C(n211), .D(n212), .Z(N298) );
  GTECH_OAI21 U227 ( .A(n192), .B(n213), .C(n214), .Z(N287) );
  GTECH_NAND3 U228 ( .A(n208), .B(n175), .C(n215), .Z(n214) );
  GTECH_NOT U229 ( .A(n176), .Z(n208) );
  GTECH_OAI21 U230 ( .A(n171), .B(n196), .C(n216), .Z(N274) );
  GTECH_NAND3 U231 ( .A(n181), .B(n191), .C(n217), .Z(n216) );
  GTECH_AND4 U232 ( .A(n215), .B(n198), .C(n169), .D(n168), .Z(N261) );
  GTECH_OAI21 U233 ( .A(n180), .B(n192), .C(n199), .Z(n198) );
  GTECH_AND2 U234 ( .A(n218), .B(n215), .Z(N248) );
  GTECH_AOI21 U235 ( .A(n169), .B(n219), .C(temp[23]), .Z(n218) );
  GTECH_NAND3 U236 ( .A(n220), .B(n199), .C(n181), .Z(n219) );
  GTECH_OAI22 U237 ( .A(n167), .B(n168), .C(n192), .D(n212), .Z(N235) );
  GTECH_NAND3 U238 ( .A(n221), .B(n220), .C(n215), .Z(n212) );
  GTECH_NOT U239 ( .A(n222), .Z(n215) );
  GTECH_NOT U240 ( .A(data_valid), .Z(n167) );
  GTECH_AND2 U241 ( .A(n156), .B(n217), .Z(N222) );
  GTECH_NOT U242 ( .A(n210), .Z(n156) );
  GTECH_NAND2 U243 ( .A(n220), .B(n186), .Z(n210) );
  GTECH_OAI21 U244 ( .A(n204), .B(n222), .C(n223), .Z(N209) );
  GTECH_NAND3 U245 ( .A(n220), .B(n188), .C(n217), .Z(n223) );
  GTECH_NOT U246 ( .A(n213), .Z(n217) );
  GTECH_NAND2 U247 ( .A(n224), .B(n225), .Z(n213) );
  GTECH_NOT U248 ( .A(n171), .Z(n224) );
  GTECH_NAND2 U249 ( .A(n157), .B(n199), .Z(n171) );
  GTECH_NOT U250 ( .A(n170), .Z(n157) );
  GTECH_NAND3 U251 ( .A(n169), .B(n168), .C(data_valid), .Z(n170) );
  GTECH_NAND2 U252 ( .A(data_valid), .B(n225), .Z(n222) );
  GTECH_NAND3 U253 ( .A(n207), .B(n190), .C(n226), .Z(n225) );
  GTECH_NOT U254 ( .A(n179), .Z(n226) );
  GTECH_NAND3 U255 ( .A(n176), .B(n204), .C(n175), .Z(n179) );
  GTECH_NAND2 U256 ( .A(temp[19]), .B(n196), .Z(n176) );
  GTECH_NAND2 U257 ( .A(n182), .B(n211), .Z(n190) );
  GTECH_NOT U258 ( .A(n227), .Z(n211) );
  GTECH_NAND2 U259 ( .A(temp[17]), .B(n186), .Z(n227) );
  GTECH_NAND3 U260 ( .A(n181), .B(n182), .C(temp[16]), .Z(n207) );
  GTECH_NOT U261 ( .A(n192), .Z(n181) );
  GTECH_NAND2 U262 ( .A(n188), .B(n186), .Z(n192) );
  GTECH_NOT U263 ( .A(temp[18]), .Z(n186) );
  GTECH_NOT U264 ( .A(temp[17]), .Z(n188) );
  GTECH_NAND2 U265 ( .A(temp[18]), .B(n182), .Z(n204) );
  GTECH_NOT U266 ( .A(n228), .Z(n182) );
  GTECH_NAND2 U267 ( .A(n175), .B(n220), .Z(n228) );
  GTECH_NOT U268 ( .A(n180), .Z(n220) );
  GTECH_NAND2 U269 ( .A(n191), .B(n196), .Z(n180) );
  GTECH_NOT U270 ( .A(temp[20]), .Z(n196) );
  GTECH_NOT U271 ( .A(temp[19]), .Z(n191) );
  GTECH_NOT U272 ( .A(n229), .Z(n175) );
  GTECH_NAND2 U273 ( .A(n221), .B(n168), .Z(n229) );
  GTECH_NOT U274 ( .A(temp[23]), .Z(n168) );
  GTECH_NOT U275 ( .A(n209), .Z(n221) );
  GTECH_NAND2 U276 ( .A(n199), .B(n169), .Z(n209) );
  GTECH_NOT U277 ( .A(temp[22]), .Z(n169) );
  GTECH_NOT U278 ( .A(temp[21]), .Z(n199) );
endmodule

