
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_XOR2 U75 ( .A(n83), .B(n84), .Z(N155) );
  GTECH_AND2 U76 ( .A(n85), .B(n86), .Z(n84) );
  GTECH_OAI22 U77 ( .A(n87), .B(n88), .C(n89), .D(n90), .Z(n83) );
  GTECH_NOT U78 ( .A(n91), .Z(n90) );
  GTECH_XOR2 U79 ( .A(n85), .B(n86), .Z(N154) );
  GTECH_NOT U80 ( .A(n92), .Z(n86) );
  GTECH_XOR2 U81 ( .A(n91), .B(n89), .Z(n92) );
  GTECH_OA21 U82 ( .A(n93), .B(n94), .C(n95), .Z(n89) );
  GTECH_OAI21 U83 ( .A(n96), .B(n97), .C(n98), .Z(n95) );
  GTECH_XOR2 U84 ( .A(n88), .B(n87), .Z(n91) );
  GTECH_OA21 U85 ( .A(n99), .B(n100), .C(n101), .Z(n87) );
  GTECH_OAI21 U86 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  GTECH_NAND2 U87 ( .A(I_b[7]), .B(I_a[7]), .Z(n88) );
  GTECH_NOT U88 ( .A(n105), .Z(n85) );
  GTECH_NAND2 U89 ( .A(n106), .B(n107), .Z(n105) );
  GTECH_XOR2 U90 ( .A(n107), .B(n106), .Z(N153) );
  GTECH_NOT U91 ( .A(n108), .Z(n106) );
  GTECH_XNOR3 U92 ( .A(n96), .B(n109), .C(n94), .Z(n108) );
  GTECH_NOT U93 ( .A(n97), .Z(n94) );
  GTECH_XNOR3 U94 ( .A(n103), .B(n102), .C(n110), .Z(n97) );
  GTECH_NOT U95 ( .A(n104), .Z(n110) );
  GTECH_OAI21 U96 ( .A(n111), .B(n112), .C(n113), .Z(n104) );
  GTECH_OAI21 U97 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_NOT U98 ( .A(n100), .Z(n102) );
  GTECH_NAND2 U99 ( .A(I_a[7]), .B(I_b[6]), .Z(n100) );
  GTECH_NOT U100 ( .A(n99), .Z(n103) );
  GTECH_NAND2 U101 ( .A(I_b[7]), .B(I_a[6]), .Z(n99) );
  GTECH_NOT U102 ( .A(n98), .Z(n109) );
  GTECH_OAI21 U103 ( .A(n117), .B(n118), .C(n119), .Z(n98) );
  GTECH_OAI21 U104 ( .A(n120), .B(n121), .C(n122), .Z(n119) );
  GTECH_NOT U105 ( .A(n93), .Z(n96) );
  GTECH_NAND2 U106 ( .A(I_a[7]), .B(n123), .Z(n93) );
  GTECH_NOT U107 ( .A(n124), .Z(n107) );
  GTECH_NAND2 U108 ( .A(n125), .B(n126), .Z(n124) );
  GTECH_XOR2 U109 ( .A(n127), .B(n128), .Z(N152) );
  GTECH_NOT U110 ( .A(n125), .Z(n128) );
  GTECH_XNOR3 U111 ( .A(n129), .B(n118), .C(n117), .Z(n125) );
  GTECH_NOT U112 ( .A(n121), .Z(n117) );
  GTECH_XOR2 U113 ( .A(n130), .B(n123), .Z(n121) );
  GTECH_OAI21 U114 ( .A(n131), .B(n132), .C(n133), .Z(n123) );
  GTECH_OAI21 U115 ( .A(n134), .B(n135), .C(n136), .Z(n133) );
  GTECH_AND2 U116 ( .A(I_a[7]), .B(I_b[5]), .Z(n130) );
  GTECH_NOT U117 ( .A(n120), .Z(n118) );
  GTECH_XNOR3 U118 ( .A(n115), .B(n114), .C(n137), .Z(n120) );
  GTECH_NOT U119 ( .A(n116), .Z(n137) );
  GTECH_OAI21 U120 ( .A(n138), .B(n139), .C(n140), .Z(n116) );
  GTECH_OAI21 U121 ( .A(n141), .B(n142), .C(n143), .Z(n140) );
  GTECH_NOT U122 ( .A(n112), .Z(n114) );
  GTECH_NAND2 U123 ( .A(I_a[6]), .B(I_b[6]), .Z(n112) );
  GTECH_NOT U124 ( .A(n111), .Z(n115) );
  GTECH_NAND2 U125 ( .A(I_b[7]), .B(I_a[5]), .Z(n111) );
  GTECH_NOT U126 ( .A(n122), .Z(n129) );
  GTECH_OAI21 U127 ( .A(n144), .B(n145), .C(n146), .Z(n122) );
  GTECH_OAI21 U128 ( .A(n147), .B(n148), .C(n149), .Z(n146) );
  GTECH_NOT U129 ( .A(n126), .Z(n127) );
  GTECH_OAI21 U130 ( .A(n150), .B(n151), .C(n152), .Z(n126) );
  GTECH_OAI21 U131 ( .A(n153), .B(n154), .C(n155), .Z(n152) );
  GTECH_XNOR3 U132 ( .A(n156), .B(n150), .C(n151), .Z(N151) );
  GTECH_NOT U133 ( .A(n153), .Z(n151) );
  GTECH_XNOR3 U134 ( .A(n157), .B(n145), .C(n144), .Z(n153) );
  GTECH_NOT U135 ( .A(n148), .Z(n144) );
  GTECH_XNOR3 U136 ( .A(n135), .B(n134), .C(n158), .Z(n148) );
  GTECH_NOT U137 ( .A(n136), .Z(n158) );
  GTECH_OAI21 U138 ( .A(n159), .B(n160), .C(n161), .Z(n136) );
  GTECH_OAI21 U139 ( .A(n162), .B(n163), .C(n164), .Z(n161) );
  GTECH_NOT U140 ( .A(n132), .Z(n134) );
  GTECH_NAND2 U141 ( .A(I_a[7]), .B(I_b[4]), .Z(n132) );
  GTECH_NOT U142 ( .A(n131), .Z(n135) );
  GTECH_NAND2 U143 ( .A(I_a[6]), .B(I_b[5]), .Z(n131) );
  GTECH_NOT U144 ( .A(n147), .Z(n145) );
  GTECH_XNOR3 U145 ( .A(n142), .B(n141), .C(n165), .Z(n147) );
  GTECH_NOT U146 ( .A(n143), .Z(n165) );
  GTECH_OAI21 U147 ( .A(n166), .B(n167), .C(n168), .Z(n143) );
  GTECH_OAI21 U148 ( .A(n169), .B(n170), .C(n171), .Z(n168) );
  GTECH_NOT U149 ( .A(n139), .Z(n141) );
  GTECH_NAND2 U150 ( .A(I_b[6]), .B(I_a[5]), .Z(n139) );
  GTECH_NOT U151 ( .A(n138), .Z(n142) );
  GTECH_NAND2 U152 ( .A(I_b[7]), .B(I_a[4]), .Z(n138) );
  GTECH_NOT U153 ( .A(n149), .Z(n157) );
  GTECH_OAI21 U154 ( .A(n172), .B(n173), .C(n174), .Z(n149) );
  GTECH_OAI21 U155 ( .A(n175), .B(n176), .C(n177), .Z(n174) );
  GTECH_NOT U156 ( .A(n154), .Z(n150) );
  GTECH_OAI22 U157 ( .A(n178), .B(n179), .C(n180), .D(n181), .Z(n154) );
  GTECH_NOT U158 ( .A(I_a[7]), .Z(n181) );
  GTECH_NOT U159 ( .A(n182), .Z(n179) );
  GTECH_NOT U160 ( .A(n155), .Z(n156) );
  GTECH_OAI2N2 U161 ( .A(n183), .B(n184), .C(n185), .D(n186), .Z(n155) );
  GTECH_OR_NOT U162 ( .A(n187), .B(n183), .Z(n186) );
  GTECH_XNOR3 U163 ( .A(n188), .B(n184), .C(n183), .Z(N150) );
  GTECH_XOR2 U164 ( .A(n182), .B(n178), .Z(n183) );
  GTECH_OA21 U165 ( .A(n189), .B(n190), .C(n191), .Z(n178) );
  GTECH_OAI21 U166 ( .A(n192), .B(n193), .C(n194), .Z(n191) );
  GTECH_XOR2 U167 ( .A(n195), .B(n180), .Z(n182) );
  GTECH_OA21 U168 ( .A(n196), .B(n197), .C(n198), .Z(n180) );
  GTECH_OAI21 U169 ( .A(n199), .B(n200), .C(n201), .Z(n198) );
  GTECH_NAND2 U170 ( .A(I_a[7]), .B(I_b[3]), .Z(n195) );
  GTECH_NOT U171 ( .A(n187), .Z(n184) );
  GTECH_XNOR3 U172 ( .A(n202), .B(n173), .C(n172), .Z(n187) );
  GTECH_NOT U173 ( .A(n176), .Z(n172) );
  GTECH_XNOR3 U174 ( .A(n163), .B(n162), .C(n203), .Z(n176) );
  GTECH_NOT U175 ( .A(n164), .Z(n203) );
  GTECH_OAI21 U176 ( .A(n204), .B(n205), .C(n206), .Z(n164) );
  GTECH_OAI21 U177 ( .A(n207), .B(n208), .C(n209), .Z(n206) );
  GTECH_NOT U178 ( .A(n160), .Z(n162) );
  GTECH_NAND2 U179 ( .A(I_a[6]), .B(I_b[4]), .Z(n160) );
  GTECH_NOT U180 ( .A(n159), .Z(n163) );
  GTECH_NAND2 U181 ( .A(I_b[5]), .B(I_a[5]), .Z(n159) );
  GTECH_NOT U182 ( .A(n175), .Z(n173) );
  GTECH_XNOR3 U183 ( .A(n170), .B(n169), .C(n210), .Z(n175) );
  GTECH_NOT U184 ( .A(n171), .Z(n210) );
  GTECH_OAI21 U185 ( .A(n211), .B(n212), .C(n213), .Z(n171) );
  GTECH_OAI21 U186 ( .A(n214), .B(n215), .C(n216), .Z(n213) );
  GTECH_NOT U187 ( .A(n167), .Z(n169) );
  GTECH_NAND2 U188 ( .A(I_b[6]), .B(I_a[4]), .Z(n167) );
  GTECH_NOT U189 ( .A(n166), .Z(n170) );
  GTECH_NAND2 U190 ( .A(I_b[7]), .B(I_a[3]), .Z(n166) );
  GTECH_NOT U191 ( .A(n177), .Z(n202) );
  GTECH_OAI21 U192 ( .A(n217), .B(n218), .C(n219), .Z(n177) );
  GTECH_OAI21 U193 ( .A(n220), .B(n221), .C(n222), .Z(n219) );
  GTECH_NOT U194 ( .A(n185), .Z(n188) );
  GTECH_OAI2N2 U195 ( .A(n223), .B(n224), .C(n225), .D(n226), .Z(n185) );
  GTECH_OR_NOT U196 ( .A(n227), .B(n223), .Z(n226) );
  GTECH_XNOR3 U197 ( .A(n228), .B(n224), .C(n223), .Z(N149) );
  GTECH_XNOR3 U198 ( .A(n192), .B(n229), .C(n190), .Z(n223) );
  GTECH_NOT U199 ( .A(n193), .Z(n190) );
  GTECH_XNOR3 U200 ( .A(n200), .B(n199), .C(n230), .Z(n193) );
  GTECH_NOT U201 ( .A(n201), .Z(n230) );
  GTECH_OAI21 U202 ( .A(n231), .B(n232), .C(n233), .Z(n201) );
  GTECH_OAI21 U203 ( .A(n234), .B(n235), .C(n236), .Z(n233) );
  GTECH_NOT U204 ( .A(n197), .Z(n199) );
  GTECH_NAND2 U205 ( .A(I_a[7]), .B(I_b[2]), .Z(n197) );
  GTECH_NOT U206 ( .A(n196), .Z(n200) );
  GTECH_NAND2 U207 ( .A(I_a[6]), .B(I_b[3]), .Z(n196) );
  GTECH_NOT U208 ( .A(n194), .Z(n229) );
  GTECH_OAI21 U209 ( .A(n237), .B(n238), .C(n239), .Z(n194) );
  GTECH_OAI21 U210 ( .A(n240), .B(n241), .C(n242), .Z(n239) );
  GTECH_NOT U211 ( .A(n189), .Z(n192) );
  GTECH_NAND2 U212 ( .A(I_a[7]), .B(n243), .Z(n189) );
  GTECH_NOT U213 ( .A(n227), .Z(n224) );
  GTECH_XNOR3 U214 ( .A(n244), .B(n218), .C(n217), .Z(n227) );
  GTECH_NOT U215 ( .A(n221), .Z(n217) );
  GTECH_XNOR3 U216 ( .A(n208), .B(n207), .C(n245), .Z(n221) );
  GTECH_NOT U217 ( .A(n209), .Z(n245) );
  GTECH_OAI21 U218 ( .A(n246), .B(n247), .C(n248), .Z(n209) );
  GTECH_OAI21 U219 ( .A(n249), .B(n250), .C(n251), .Z(n248) );
  GTECH_NOT U220 ( .A(n205), .Z(n207) );
  GTECH_NAND2 U221 ( .A(I_a[5]), .B(I_b[4]), .Z(n205) );
  GTECH_NOT U222 ( .A(n204), .Z(n208) );
  GTECH_NAND2 U223 ( .A(I_b[5]), .B(I_a[4]), .Z(n204) );
  GTECH_NOT U224 ( .A(n220), .Z(n218) );
  GTECH_XNOR3 U225 ( .A(n215), .B(n214), .C(n252), .Z(n220) );
  GTECH_NOT U226 ( .A(n216), .Z(n252) );
  GTECH_OAI21 U227 ( .A(n253), .B(n254), .C(n255), .Z(n216) );
  GTECH_NOT U228 ( .A(n212), .Z(n214) );
  GTECH_NAND2 U229 ( .A(I_b[6]), .B(I_a[3]), .Z(n212) );
  GTECH_NOT U230 ( .A(n211), .Z(n215) );
  GTECH_NAND2 U231 ( .A(I_b[7]), .B(I_a[2]), .Z(n211) );
  GTECH_NOT U232 ( .A(n222), .Z(n244) );
  GTECH_OAI21 U233 ( .A(n256), .B(n257), .C(n258), .Z(n222) );
  GTECH_OAI21 U234 ( .A(n259), .B(n260), .C(n261), .Z(n258) );
  GTECH_NOT U235 ( .A(n225), .Z(n228) );
  GTECH_OAI2N2 U236 ( .A(n262), .B(n263), .C(n264), .D(n265), .Z(n225) );
  GTECH_OR_NOT U237 ( .A(n266), .B(n262), .Z(n265) );
  GTECH_XNOR3 U238 ( .A(n267), .B(n263), .C(n262), .Z(N148) );
  GTECH_XNOR3 U239 ( .A(n268), .B(n257), .C(n260), .Z(n262) );
  GTECH_NOT U240 ( .A(n256), .Z(n260) );
  GTECH_XNOR3 U241 ( .A(n269), .B(n270), .C(n271), .Z(n256) );
  GTECH_NOT U242 ( .A(n255), .Z(n271) );
  GTECH_NAND3 U243 ( .A(I_b[6]), .B(I_a[1]), .C(n272), .Z(n255) );
  GTECH_NOT U244 ( .A(n254), .Z(n270) );
  GTECH_NAND2 U245 ( .A(I_b[6]), .B(I_a[2]), .Z(n254) );
  GTECH_NOT U246 ( .A(n253), .Z(n269) );
  GTECH_NAND2 U247 ( .A(I_b[7]), .B(I_a[1]), .Z(n253) );
  GTECH_NOT U248 ( .A(n259), .Z(n257) );
  GTECH_XNOR3 U249 ( .A(n250), .B(n249), .C(n273), .Z(n259) );
  GTECH_NOT U250 ( .A(n251), .Z(n273) );
  GTECH_OAI21 U251 ( .A(n274), .B(n275), .C(n276), .Z(n251) );
  GTECH_OAI21 U252 ( .A(n277), .B(n278), .C(n279), .Z(n276) );
  GTECH_NOT U253 ( .A(n247), .Z(n249) );
  GTECH_NAND2 U254 ( .A(I_b[4]), .B(I_a[4]), .Z(n247) );
  GTECH_NOT U255 ( .A(n246), .Z(n250) );
  GTECH_NAND2 U256 ( .A(I_b[5]), .B(I_a[3]), .Z(n246) );
  GTECH_NOT U257 ( .A(n261), .Z(n268) );
  GTECH_OAI21 U258 ( .A(n280), .B(n281), .C(n282), .Z(n261) );
  GTECH_OAI21 U259 ( .A(n283), .B(n284), .C(n285), .Z(n282) );
  GTECH_NOT U260 ( .A(n266), .Z(n263) );
  GTECH_XNOR3 U261 ( .A(n286), .B(n238), .C(n237), .Z(n266) );
  GTECH_NOT U262 ( .A(n241), .Z(n237) );
  GTECH_XOR2 U263 ( .A(n287), .B(n243), .Z(n241) );
  GTECH_OAI21 U264 ( .A(n288), .B(n289), .C(n290), .Z(n243) );
  GTECH_OAI21 U265 ( .A(n291), .B(n292), .C(n293), .Z(n290) );
  GTECH_AND2 U266 ( .A(I_a[7]), .B(I_b[1]), .Z(n287) );
  GTECH_NOT U267 ( .A(n240), .Z(n238) );
  GTECH_XNOR3 U268 ( .A(n235), .B(n234), .C(n294), .Z(n240) );
  GTECH_NOT U269 ( .A(n236), .Z(n294) );
  GTECH_OAI21 U270 ( .A(n295), .B(n296), .C(n297), .Z(n236) );
  GTECH_OAI21 U271 ( .A(n298), .B(n299), .C(n300), .Z(n297) );
  GTECH_NOT U272 ( .A(n232), .Z(n234) );
  GTECH_NAND2 U273 ( .A(I_a[6]), .B(I_b[2]), .Z(n232) );
  GTECH_NOT U274 ( .A(n231), .Z(n235) );
  GTECH_NAND2 U275 ( .A(I_a[5]), .B(I_b[3]), .Z(n231) );
  GTECH_NOT U276 ( .A(n242), .Z(n286) );
  GTECH_OAI21 U277 ( .A(n301), .B(n302), .C(n303), .Z(n242) );
  GTECH_OAI21 U278 ( .A(n304), .B(n305), .C(n306), .Z(n303) );
  GTECH_NOT U279 ( .A(n264), .Z(n267) );
  GTECH_OAI21 U280 ( .A(n307), .B(n308), .C(n309), .Z(n264) );
  GTECH_OAI21 U281 ( .A(n310), .B(n311), .C(n312), .Z(n309) );
  GTECH_XNOR3 U282 ( .A(n313), .B(n308), .C(n307), .Z(N147) );
  GTECH_NOT U283 ( .A(n311), .Z(n307) );
  GTECH_XNOR3 U284 ( .A(n285), .B(n281), .C(n284), .Z(n311) );
  GTECH_NOT U285 ( .A(n280), .Z(n284) );
  GTECH_XOR2 U286 ( .A(n314), .B(n272), .Z(n280) );
  GTECH_NOT U287 ( .A(n315), .Z(n272) );
  GTECH_NAND2 U288 ( .A(I_b[7]), .B(I_a[0]), .Z(n315) );
  GTECH_NAND2 U289 ( .A(I_b[6]), .B(I_a[1]), .Z(n314) );
  GTECH_NOT U290 ( .A(n283), .Z(n281) );
  GTECH_XNOR3 U291 ( .A(n278), .B(n277), .C(n316), .Z(n283) );
  GTECH_NOT U292 ( .A(n279), .Z(n316) );
  GTECH_OAI21 U293 ( .A(n317), .B(n318), .C(n319), .Z(n279) );
  GTECH_NOT U294 ( .A(n275), .Z(n277) );
  GTECH_NAND2 U295 ( .A(I_b[4]), .B(I_a[3]), .Z(n275) );
  GTECH_NOT U296 ( .A(n274), .Z(n278) );
  GTECH_NAND2 U297 ( .A(I_b[5]), .B(I_a[2]), .Z(n274) );
  GTECH_NOT U298 ( .A(n320), .Z(n285) );
  GTECH_NOT U299 ( .A(n310), .Z(n308) );
  GTECH_XNOR3 U300 ( .A(n321), .B(n302), .C(n301), .Z(n310) );
  GTECH_NOT U301 ( .A(n305), .Z(n301) );
  GTECH_XNOR3 U302 ( .A(n299), .B(n298), .C(n322), .Z(n305) );
  GTECH_NOT U303 ( .A(n300), .Z(n322) );
  GTECH_OAI21 U304 ( .A(n323), .B(n324), .C(n325), .Z(n300) );
  GTECH_OAI21 U305 ( .A(n326), .B(n327), .C(n328), .Z(n325) );
  GTECH_NOT U306 ( .A(n296), .Z(n298) );
  GTECH_NAND2 U307 ( .A(I_a[5]), .B(I_b[2]), .Z(n296) );
  GTECH_NOT U308 ( .A(n295), .Z(n299) );
  GTECH_NAND2 U309 ( .A(I_a[4]), .B(I_b[3]), .Z(n295) );
  GTECH_NOT U310 ( .A(n304), .Z(n302) );
  GTECH_XNOR3 U311 ( .A(n292), .B(n291), .C(n329), .Z(n304) );
  GTECH_NOT U312 ( .A(n293), .Z(n329) );
  GTECH_OAI21 U313 ( .A(n330), .B(n331), .C(n332), .Z(n293) );
  GTECH_OAI21 U314 ( .A(n333), .B(n334), .C(n335), .Z(n332) );
  GTECH_NOT U315 ( .A(n289), .Z(n291) );
  GTECH_NAND2 U316 ( .A(I_a[7]), .B(I_b[0]), .Z(n289) );
  GTECH_NOT U317 ( .A(n288), .Z(n292) );
  GTECH_NAND2 U318 ( .A(I_a[6]), .B(I_b[1]), .Z(n288) );
  GTECH_NOT U319 ( .A(n306), .Z(n321) );
  GTECH_OAI21 U320 ( .A(n336), .B(n337), .C(n338), .Z(n306) );
  GTECH_OAI21 U321 ( .A(n339), .B(n340), .C(n341), .Z(n338) );
  GTECH_NOT U322 ( .A(n312), .Z(n313) );
  GTECH_OAI21 U323 ( .A(n342), .B(n343), .C(n344), .Z(n312) );
  GTECH_OAI21 U324 ( .A(n345), .B(n346), .C(n347), .Z(n344) );
  GTECH_NOT U325 ( .A(n346), .Z(n342) );
  GTECH_XNOR3 U326 ( .A(n345), .B(n348), .C(n346), .Z(N146) );
  GTECH_XNOR3 U327 ( .A(n349), .B(n337), .C(n336), .Z(n346) );
  GTECH_NOT U328 ( .A(n340), .Z(n336) );
  GTECH_XNOR3 U329 ( .A(n327), .B(n326), .C(n350), .Z(n340) );
  GTECH_NOT U330 ( .A(n328), .Z(n350) );
  GTECH_OAI21 U331 ( .A(n351), .B(n352), .C(n353), .Z(n328) );
  GTECH_OAI21 U332 ( .A(n354), .B(n355), .C(n356), .Z(n353) );
  GTECH_NOT U333 ( .A(n324), .Z(n326) );
  GTECH_NAND2 U334 ( .A(I_a[4]), .B(I_b[2]), .Z(n324) );
  GTECH_NOT U335 ( .A(n323), .Z(n327) );
  GTECH_NAND2 U336 ( .A(I_a[3]), .B(I_b[3]), .Z(n323) );
  GTECH_NOT U337 ( .A(n339), .Z(n337) );
  GTECH_XNOR3 U338 ( .A(n334), .B(n333), .C(n357), .Z(n339) );
  GTECH_NOT U339 ( .A(n335), .Z(n357) );
  GTECH_OAI21 U340 ( .A(n358), .B(n359), .C(n360), .Z(n335) );
  GTECH_OAI21 U341 ( .A(n361), .B(n362), .C(n363), .Z(n360) );
  GTECH_NOT U342 ( .A(n331), .Z(n333) );
  GTECH_NAND2 U343 ( .A(I_a[6]), .B(I_b[0]), .Z(n331) );
  GTECH_NOT U344 ( .A(n330), .Z(n334) );
  GTECH_NAND2 U345 ( .A(I_a[5]), .B(I_b[1]), .Z(n330) );
  GTECH_NOT U346 ( .A(n341), .Z(n349) );
  GTECH_OAI21 U347 ( .A(n364), .B(n365), .C(n366), .Z(n341) );
  GTECH_OAI21 U348 ( .A(n367), .B(n368), .C(n369), .Z(n366) );
  GTECH_NOT U349 ( .A(n347), .Z(n348) );
  GTECH_OAI21 U350 ( .A(n370), .B(n371), .C(n372), .Z(n347) );
  GTECH_OAI21 U351 ( .A(n373), .B(n374), .C(n375), .Z(n372) );
  GTECH_NOT U352 ( .A(n343), .Z(n345) );
  GTECH_NAND2 U353 ( .A(n320), .B(n376), .Z(n343) );
  GTECH_NAND2 U354 ( .A(n377), .B(n378), .Z(n376) );
  GTECH_NAND2 U355 ( .A(I_a[0]), .B(I_b[6]), .Z(n378) );
  GTECH_NAND3 U356 ( .A(I_a[0]), .B(n379), .C(I_b[6]), .Z(n320) );
  GTECH_NOT U357 ( .A(n377), .Z(n379) );
  GTECH_XNOR3 U358 ( .A(n380), .B(n381), .C(n382), .Z(n377) );
  GTECH_NOT U359 ( .A(n319), .Z(n382) );
  GTECH_NAND3 U360 ( .A(I_b[4]), .B(I_a[1]), .C(n383), .Z(n319) );
  GTECH_NOT U361 ( .A(n318), .Z(n381) );
  GTECH_NAND2 U362 ( .A(I_b[4]), .B(I_a[2]), .Z(n318) );
  GTECH_NOT U363 ( .A(n317), .Z(n380) );
  GTECH_NAND2 U364 ( .A(I_b[5]), .B(I_a[1]), .Z(n317) );
  GTECH_XNOR3 U365 ( .A(n375), .B(n371), .C(n374), .Z(N145) );
  GTECH_NOT U366 ( .A(n370), .Z(n374) );
  GTECH_XOR2 U367 ( .A(n384), .B(n383), .Z(n370) );
  GTECH_NOT U368 ( .A(n385), .Z(n383) );
  GTECH_NAND2 U369 ( .A(I_b[5]), .B(I_a[0]), .Z(n385) );
  GTECH_NAND2 U370 ( .A(I_b[4]), .B(I_a[1]), .Z(n384) );
  GTECH_NOT U371 ( .A(n373), .Z(n371) );
  GTECH_XNOR3 U372 ( .A(n386), .B(n365), .C(n364), .Z(n373) );
  GTECH_NOT U373 ( .A(n368), .Z(n364) );
  GTECH_XNOR3 U374 ( .A(n362), .B(n361), .C(n387), .Z(n368) );
  GTECH_NOT U375 ( .A(n363), .Z(n387) );
  GTECH_OAI21 U376 ( .A(n388), .B(n389), .C(n390), .Z(n363) );
  GTECH_OAI21 U377 ( .A(n391), .B(n392), .C(n393), .Z(n390) );
  GTECH_NOT U378 ( .A(n359), .Z(n361) );
  GTECH_NAND2 U379 ( .A(I_a[5]), .B(I_b[0]), .Z(n359) );
  GTECH_NOT U380 ( .A(n358), .Z(n362) );
  GTECH_NAND2 U381 ( .A(I_a[4]), .B(I_b[1]), .Z(n358) );
  GTECH_NOT U382 ( .A(n367), .Z(n365) );
  GTECH_XNOR3 U383 ( .A(n355), .B(n354), .C(n394), .Z(n367) );
  GTECH_NOT U384 ( .A(n356), .Z(n394) );
  GTECH_OAI21 U385 ( .A(n395), .B(n396), .C(n397), .Z(n356) );
  GTECH_NOT U386 ( .A(n352), .Z(n354) );
  GTECH_NAND2 U387 ( .A(I_a[3]), .B(I_b[2]), .Z(n352) );
  GTECH_NOT U388 ( .A(n351), .Z(n355) );
  GTECH_NAND2 U389 ( .A(I_a[2]), .B(I_b[3]), .Z(n351) );
  GTECH_NOT U390 ( .A(n369), .Z(n386) );
  GTECH_OAI21 U391 ( .A(n398), .B(n399), .C(n400), .Z(n369) );
  GTECH_OAI21 U392 ( .A(n401), .B(n402), .C(n403), .Z(n400) );
  GTECH_NOT U393 ( .A(n404), .Z(n375) );
  GTECH_NAND3 U394 ( .A(I_a[0]), .B(n405), .C(I_b[4]), .Z(n404) );
  GTECH_XOR2 U395 ( .A(n406), .B(n405), .Z(N144) );
  GTECH_NOT U396 ( .A(n407), .Z(n405) );
  GTECH_XNOR3 U397 ( .A(n408), .B(n399), .C(n402), .Z(n407) );
  GTECH_NOT U398 ( .A(n398), .Z(n402) );
  GTECH_XNOR3 U399 ( .A(n409), .B(n410), .C(n411), .Z(n398) );
  GTECH_NOT U400 ( .A(n397), .Z(n411) );
  GTECH_NAND3 U401 ( .A(I_a[1]), .B(n412), .C(I_b[2]), .Z(n397) );
  GTECH_NOT U402 ( .A(n396), .Z(n410) );
  GTECH_NAND2 U403 ( .A(I_a[2]), .B(I_b[2]), .Z(n396) );
  GTECH_NOT U404 ( .A(n395), .Z(n409) );
  GTECH_NAND2 U405 ( .A(I_a[1]), .B(I_b[3]), .Z(n395) );
  GTECH_NOT U406 ( .A(n401), .Z(n399) );
  GTECH_XNOR3 U407 ( .A(n392), .B(n391), .C(n413), .Z(n401) );
  GTECH_NOT U408 ( .A(n393), .Z(n413) );
  GTECH_OAI21 U409 ( .A(n414), .B(n415), .C(n416), .Z(n393) );
  GTECH_OAI21 U410 ( .A(n417), .B(n418), .C(n419), .Z(n416) );
  GTECH_NOT U411 ( .A(n389), .Z(n391) );
  GTECH_NAND2 U412 ( .A(I_a[4]), .B(I_b[0]), .Z(n389) );
  GTECH_NOT U413 ( .A(n388), .Z(n392) );
  GTECH_NAND2 U414 ( .A(I_a[3]), .B(I_b[1]), .Z(n388) );
  GTECH_NOT U415 ( .A(n403), .Z(n408) );
  GTECH_OAI21 U416 ( .A(n420), .B(n421), .C(n422), .Z(n403) );
  GTECH_OAI21 U417 ( .A(n423), .B(n424), .C(n425), .Z(n422) );
  GTECH_AND2 U418 ( .A(I_b[4]), .B(I_a[0]), .Z(n406) );
  GTECH_XNOR3 U419 ( .A(n425), .B(n421), .C(n424), .Z(N143) );
  GTECH_NOT U420 ( .A(n420), .Z(n424) );
  GTECH_XOR2 U421 ( .A(n426), .B(n412), .Z(n420) );
  GTECH_NOT U422 ( .A(n427), .Z(n412) );
  GTECH_NAND2 U423 ( .A(I_b[3]), .B(I_a[0]), .Z(n427) );
  GTECH_NAND2 U424 ( .A(I_b[2]), .B(I_a[1]), .Z(n426) );
  GTECH_NOT U425 ( .A(n423), .Z(n421) );
  GTECH_XNOR3 U426 ( .A(n418), .B(n417), .C(n428), .Z(n423) );
  GTECH_NOT U427 ( .A(n419), .Z(n428) );
  GTECH_OAI21 U428 ( .A(n429), .B(n430), .C(n431), .Z(n419) );
  GTECH_NOT U429 ( .A(n415), .Z(n417) );
  GTECH_NAND2 U430 ( .A(I_a[3]), .B(I_b[0]), .Z(n415) );
  GTECH_NOT U431 ( .A(n414), .Z(n418) );
  GTECH_NAND2 U432 ( .A(I_b[1]), .B(I_a[2]), .Z(n414) );
  GTECH_NOT U433 ( .A(n432), .Z(n425) );
  GTECH_NAND3 U434 ( .A(I_a[0]), .B(n433), .C(I_b[2]), .Z(n432) );
  GTECH_XOR2 U435 ( .A(n434), .B(n433), .Z(N142) );
  GTECH_NOT U436 ( .A(n435), .Z(n433) );
  GTECH_XNOR3 U437 ( .A(n436), .B(n437), .C(n438), .Z(n435) );
  GTECH_NOT U438 ( .A(n431), .Z(n438) );
  GTECH_NAND3 U439 ( .A(n439), .B(I_a[1]), .C(I_b[0]), .Z(n431) );
  GTECH_NOT U440 ( .A(n430), .Z(n437) );
  GTECH_NAND2 U441 ( .A(I_b[0]), .B(I_a[2]), .Z(n430) );
  GTECH_NOT U442 ( .A(n429), .Z(n436) );
  GTECH_NAND2 U443 ( .A(I_b[1]), .B(I_a[1]), .Z(n429) );
  GTECH_AND2 U444 ( .A(I_b[2]), .B(I_a[0]), .Z(n434) );
  GTECH_XOR2 U445 ( .A(n439), .B(n440), .Z(N141) );
  GTECH_AND2 U446 ( .A(I_b[0]), .B(I_a[1]), .Z(n440) );
  GTECH_NOT U447 ( .A(n441), .Z(n439) );
  GTECH_NAND2 U448 ( .A(I_b[1]), .B(I_a[0]), .Z(n441) );
  GTECH_AND2 U449 ( .A(I_b[0]), .B(I_a[0]), .Z(N140) );
endmodule

