
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_XNOR2 U75 ( .A(n83), .B(n84), .Z(N155) );
  GTECH_OA22 U76 ( .A(n85), .B(n86), .C(n87), .D(n88), .Z(n84) );
  GTECH_AND_NOT U77 ( .A(n89), .B(n90), .Z(n83) );
  GTECH_XNOR2 U78 ( .A(n89), .B(n90), .Z(N154) );
  GTECH_XNOR2 U79 ( .A(n88), .B(n87), .Z(n90) );
  GTECH_NOT U80 ( .A(n91), .Z(n87) );
  GTECH_XNOR2 U81 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U82 ( .A(n85), .Z(n92) );
  GTECH_NAND2 U83 ( .A(I_b[7]), .B(I_a[7]), .Z(n85) );
  GTECH_OA21 U84 ( .A(n93), .B(n94), .C(n95), .Z(n86) );
  GTECH_OAI21 U85 ( .A(n96), .B(n97), .C(n98), .Z(n95) );
  GTECH_AND2 U86 ( .A(n99), .B(n100), .Z(n88) );
  GTECH_OR_NOT U87 ( .A(n101), .B(n102), .Z(n100) );
  GTECH_OAI21 U88 ( .A(n103), .B(n102), .C(n104), .Z(n99) );
  GTECH_NOT U89 ( .A(n105), .Z(n89) );
  GTECH_NAND2 U90 ( .A(n106), .B(n107), .Z(n105) );
  GTECH_NOT U91 ( .A(n108), .Z(n106) );
  GTECH_XNOR2 U92 ( .A(n107), .B(n108), .Z(N153) );
  GTECH_XOR3 U93 ( .A(n103), .B(n109), .C(n102), .Z(n108) );
  GTECH_XOR3 U94 ( .A(n97), .B(n96), .C(n98), .Z(n102) );
  GTECH_OAI21 U95 ( .A(n110), .B(n111), .C(n112), .Z(n98) );
  GTECH_OAI21 U96 ( .A(n113), .B(n114), .C(n115), .Z(n112) );
  GTECH_NOT U97 ( .A(n94), .Z(n96) );
  GTECH_NAND2 U98 ( .A(I_a[7]), .B(I_b[6]), .Z(n94) );
  GTECH_NOT U99 ( .A(n93), .Z(n97) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n93) );
  GTECH_NOT U101 ( .A(n104), .Z(n109) );
  GTECH_AO22 U102 ( .A(n116), .B(n117), .C(n118), .D(n119), .Z(n104) );
  GTECH_OR2 U103 ( .A(n119), .B(n118), .Z(n117) );
  GTECH_NOT U104 ( .A(n101), .Z(n103) );
  GTECH_NAND2 U105 ( .A(I_a[7]), .B(n120), .Z(n101) );
  GTECH_NOT U106 ( .A(n121), .Z(n107) );
  GTECH_NAND2 U107 ( .A(n122), .B(n123), .Z(n121) );
  GTECH_XNOR2 U108 ( .A(n124), .B(n122), .Z(N152) );
  GTECH_XOR3 U109 ( .A(n125), .B(n126), .C(n118), .Z(n122) );
  GTECH_XNOR2 U110 ( .A(n120), .B(n127), .Z(n118) );
  GTECH_NAND2 U111 ( .A(I_a[7]), .B(I_b[5]), .Z(n127) );
  GTECH_OAI21 U112 ( .A(n128), .B(n129), .C(n130), .Z(n120) );
  GTECH_OAI21 U113 ( .A(n131), .B(n132), .C(n133), .Z(n130) );
  GTECH_NOT U114 ( .A(n119), .Z(n126) );
  GTECH_XOR3 U115 ( .A(n114), .B(n113), .C(n115), .Z(n119) );
  GTECH_OAI21 U116 ( .A(n134), .B(n135), .C(n136), .Z(n115) );
  GTECH_OAI21 U117 ( .A(n137), .B(n138), .C(n139), .Z(n136) );
  GTECH_NOT U118 ( .A(n111), .Z(n113) );
  GTECH_NAND2 U119 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_NOT U120 ( .A(n110), .Z(n114) );
  GTECH_NAND2 U121 ( .A(I_b[7]), .B(I_a[5]), .Z(n110) );
  GTECH_NOT U122 ( .A(n116), .Z(n125) );
  GTECH_AO22 U123 ( .A(n140), .B(n141), .C(n142), .D(n143), .Z(n116) );
  GTECH_OR2 U124 ( .A(n143), .B(n142), .Z(n141) );
  GTECH_NOT U125 ( .A(n123), .Z(n124) );
  GTECH_AO22 U126 ( .A(n144), .B(n145), .C(n146), .D(n147), .Z(n123) );
  GTECH_OR2 U127 ( .A(n146), .B(n147), .Z(n145) );
  GTECH_XOR3 U128 ( .A(n148), .B(n149), .C(n146), .Z(N151) );
  GTECH_XOR3 U129 ( .A(n150), .B(n151), .C(n142), .Z(n146) );
  GTECH_XOR3 U130 ( .A(n132), .B(n131), .C(n133), .Z(n142) );
  GTECH_OAI21 U131 ( .A(n152), .B(n153), .C(n154), .Z(n133) );
  GTECH_OAI21 U132 ( .A(n155), .B(n156), .C(n157), .Z(n154) );
  GTECH_NOT U133 ( .A(n129), .Z(n131) );
  GTECH_NAND2 U134 ( .A(I_a[7]), .B(I_b[4]), .Z(n129) );
  GTECH_NOT U135 ( .A(n128), .Z(n132) );
  GTECH_NAND2 U136 ( .A(I_a[6]), .B(I_b[5]), .Z(n128) );
  GTECH_NOT U137 ( .A(n143), .Z(n151) );
  GTECH_XOR3 U138 ( .A(n138), .B(n137), .C(n139), .Z(n143) );
  GTECH_OAI21 U139 ( .A(n158), .B(n159), .C(n160), .Z(n139) );
  GTECH_OAI21 U140 ( .A(n161), .B(n162), .C(n163), .Z(n160) );
  GTECH_NOT U141 ( .A(n135), .Z(n137) );
  GTECH_NAND2 U142 ( .A(I_b[6]), .B(I_a[5]), .Z(n135) );
  GTECH_NOT U143 ( .A(n134), .Z(n138) );
  GTECH_NAND2 U144 ( .A(I_b[7]), .B(I_a[4]), .Z(n134) );
  GTECH_NOT U145 ( .A(n140), .Z(n150) );
  GTECH_AO22 U146 ( .A(n164), .B(n165), .C(n166), .D(n167), .Z(n140) );
  GTECH_OR2 U147 ( .A(n167), .B(n166), .Z(n165) );
  GTECH_NOT U148 ( .A(n147), .Z(n149) );
  GTECH_OAI22 U149 ( .A(n168), .B(n169), .C(n170), .D(n171), .Z(n147) );
  GTECH_NOT U150 ( .A(I_a[7]), .Z(n171) );
  GTECH_NOT U151 ( .A(n144), .Z(n148) );
  GTECH_OAI21 U152 ( .A(n172), .B(n173), .C(n174), .Z(n144) );
  GTECH_OAI21 U153 ( .A(n175), .B(n176), .C(n177), .Z(n174) );
  GTECH_XOR3 U154 ( .A(n178), .B(n173), .C(n176), .Z(N150) );
  GTECH_NOT U155 ( .A(n172), .Z(n176) );
  GTECH_XNOR2 U156 ( .A(n168), .B(n169), .Z(n172) );
  GTECH_XNOR2 U157 ( .A(n170), .B(n179), .Z(n169) );
  GTECH_NAND2 U158 ( .A(I_a[7]), .B(I_b[3]), .Z(n179) );
  GTECH_OA21 U159 ( .A(n180), .B(n181), .C(n182), .Z(n170) );
  GTECH_OAI21 U160 ( .A(n183), .B(n184), .C(n185), .Z(n182) );
  GTECH_AND2 U161 ( .A(n186), .B(n187), .Z(n168) );
  GTECH_OR_NOT U162 ( .A(n188), .B(n189), .Z(n187) );
  GTECH_OAI21 U163 ( .A(n190), .B(n189), .C(n191), .Z(n186) );
  GTECH_NOT U164 ( .A(n175), .Z(n173) );
  GTECH_XOR3 U165 ( .A(n192), .B(n193), .C(n166), .Z(n175) );
  GTECH_XOR3 U166 ( .A(n156), .B(n155), .C(n157), .Z(n166) );
  GTECH_OAI21 U167 ( .A(n194), .B(n195), .C(n196), .Z(n157) );
  GTECH_OAI21 U168 ( .A(n197), .B(n198), .C(n199), .Z(n196) );
  GTECH_NOT U169 ( .A(n153), .Z(n155) );
  GTECH_NAND2 U170 ( .A(I_a[6]), .B(I_b[4]), .Z(n153) );
  GTECH_NOT U171 ( .A(n152), .Z(n156) );
  GTECH_NAND2 U172 ( .A(I_b[5]), .B(I_a[5]), .Z(n152) );
  GTECH_NOT U173 ( .A(n167), .Z(n193) );
  GTECH_XOR3 U174 ( .A(n162), .B(n161), .C(n163), .Z(n167) );
  GTECH_OAI21 U175 ( .A(n200), .B(n201), .C(n202), .Z(n163) );
  GTECH_OAI21 U176 ( .A(n203), .B(n204), .C(n205), .Z(n202) );
  GTECH_NOT U177 ( .A(n159), .Z(n161) );
  GTECH_NAND2 U178 ( .A(I_b[6]), .B(I_a[4]), .Z(n159) );
  GTECH_NOT U179 ( .A(n158), .Z(n162) );
  GTECH_NAND2 U180 ( .A(I_b[7]), .B(I_a[3]), .Z(n158) );
  GTECH_NOT U181 ( .A(n164), .Z(n192) );
  GTECH_AO22 U182 ( .A(n206), .B(n207), .C(n208), .D(n209), .Z(n164) );
  GTECH_OR2 U183 ( .A(n209), .B(n208), .Z(n207) );
  GTECH_NOT U184 ( .A(n177), .Z(n178) );
  GTECH_OAI21 U185 ( .A(n210), .B(n211), .C(n212), .Z(n177) );
  GTECH_OAI21 U186 ( .A(n213), .B(n214), .C(n215), .Z(n212) );
  GTECH_XOR3 U187 ( .A(n216), .B(n211), .C(n214), .Z(N149) );
  GTECH_NOT U188 ( .A(n210), .Z(n214) );
  GTECH_XOR3 U189 ( .A(n190), .B(n217), .C(n189), .Z(n210) );
  GTECH_XOR3 U190 ( .A(n184), .B(n183), .C(n185), .Z(n189) );
  GTECH_OAI21 U191 ( .A(n218), .B(n219), .C(n220), .Z(n185) );
  GTECH_OAI21 U192 ( .A(n221), .B(n222), .C(n223), .Z(n220) );
  GTECH_NOT U193 ( .A(n181), .Z(n183) );
  GTECH_NAND2 U194 ( .A(I_a[7]), .B(I_b[2]), .Z(n181) );
  GTECH_NOT U195 ( .A(n180), .Z(n184) );
  GTECH_NAND2 U196 ( .A(I_a[6]), .B(I_b[3]), .Z(n180) );
  GTECH_NOT U197 ( .A(n191), .Z(n217) );
  GTECH_AO22 U198 ( .A(n224), .B(n225), .C(n226), .D(n227), .Z(n191) );
  GTECH_OR2 U199 ( .A(n227), .B(n226), .Z(n225) );
  GTECH_NOT U200 ( .A(n188), .Z(n190) );
  GTECH_NAND2 U201 ( .A(I_a[7]), .B(n228), .Z(n188) );
  GTECH_NOT U202 ( .A(n213), .Z(n211) );
  GTECH_XOR3 U203 ( .A(n229), .B(n230), .C(n208), .Z(n213) );
  GTECH_XOR3 U204 ( .A(n198), .B(n197), .C(n199), .Z(n208) );
  GTECH_OAI21 U205 ( .A(n231), .B(n232), .C(n233), .Z(n199) );
  GTECH_OAI21 U206 ( .A(n234), .B(n235), .C(n236), .Z(n233) );
  GTECH_NOT U207 ( .A(n195), .Z(n197) );
  GTECH_NAND2 U208 ( .A(I_a[5]), .B(I_b[4]), .Z(n195) );
  GTECH_NOT U209 ( .A(n194), .Z(n198) );
  GTECH_NAND2 U210 ( .A(I_b[5]), .B(I_a[4]), .Z(n194) );
  GTECH_NOT U211 ( .A(n209), .Z(n230) );
  GTECH_XOR3 U212 ( .A(n204), .B(n203), .C(n205), .Z(n209) );
  GTECH_OAI21 U213 ( .A(n237), .B(n238), .C(n239), .Z(n205) );
  GTECH_NOT U214 ( .A(n201), .Z(n203) );
  GTECH_NAND2 U215 ( .A(I_b[6]), .B(I_a[3]), .Z(n201) );
  GTECH_NOT U216 ( .A(n200), .Z(n204) );
  GTECH_NAND2 U217 ( .A(I_b[7]), .B(I_a[2]), .Z(n200) );
  GTECH_NOT U218 ( .A(n206), .Z(n229) );
  GTECH_OAI2N2 U219 ( .A(n240), .B(n241), .C(n242), .D(n243), .Z(n206) );
  GTECH_OR_NOT U220 ( .A(n244), .B(n240), .Z(n243) );
  GTECH_NOT U221 ( .A(n215), .Z(n216) );
  GTECH_OAI21 U222 ( .A(n245), .B(n246), .C(n247), .Z(n215) );
  GTECH_OAI21 U223 ( .A(n248), .B(n249), .C(n250), .Z(n247) );
  GTECH_XOR3 U224 ( .A(n251), .B(n246), .C(n249), .Z(N148) );
  GTECH_NOT U225 ( .A(n245), .Z(n249) );
  GTECH_XOR3 U226 ( .A(n252), .B(n241), .C(n240), .Z(n245) );
  GTECH_XOR3 U227 ( .A(n253), .B(n254), .C(n239), .Z(n240) );
  GTECH_NAND3 U228 ( .A(I_b[7]), .B(I_a[0]), .C(n255), .Z(n239) );
  GTECH_NOT U229 ( .A(n238), .Z(n254) );
  GTECH_NAND2 U230 ( .A(I_b[6]), .B(I_a[2]), .Z(n238) );
  GTECH_NOT U231 ( .A(n237), .Z(n253) );
  GTECH_NAND2 U232 ( .A(I_b[7]), .B(I_a[1]), .Z(n237) );
  GTECH_NOT U233 ( .A(n244), .Z(n241) );
  GTECH_XOR3 U234 ( .A(n235), .B(n234), .C(n236), .Z(n244) );
  GTECH_OAI21 U235 ( .A(n256), .B(n257), .C(n258), .Z(n236) );
  GTECH_OAI21 U236 ( .A(n259), .B(n260), .C(n261), .Z(n258) );
  GTECH_NOT U237 ( .A(n232), .Z(n234) );
  GTECH_NAND2 U238 ( .A(I_b[4]), .B(I_a[4]), .Z(n232) );
  GTECH_NOT U239 ( .A(n231), .Z(n235) );
  GTECH_NAND2 U240 ( .A(I_b[5]), .B(I_a[3]), .Z(n231) );
  GTECH_NOT U241 ( .A(n242), .Z(n252) );
  GTECH_OAI22 U242 ( .A(n262), .B(n263), .C(n264), .D(n265), .Z(n242) );
  GTECH_AND_NOT U243 ( .A(n264), .B(n266), .Z(n262) );
  GTECH_NOT U244 ( .A(n248), .Z(n246) );
  GTECH_XOR3 U245 ( .A(n267), .B(n268), .C(n226), .Z(n248) );
  GTECH_XNOR2 U246 ( .A(n228), .B(n269), .Z(n226) );
  GTECH_NAND2 U247 ( .A(I_a[7]), .B(I_b[1]), .Z(n269) );
  GTECH_OAI21 U248 ( .A(n270), .B(n271), .C(n272), .Z(n228) );
  GTECH_AO21 U249 ( .A(n270), .B(n271), .C(n273), .Z(n272) );
  GTECH_NOT U250 ( .A(n227), .Z(n268) );
  GTECH_XOR3 U251 ( .A(n222), .B(n221), .C(n223), .Z(n227) );
  GTECH_OAI21 U252 ( .A(n274), .B(n275), .C(n276), .Z(n223) );
  GTECH_OAI21 U253 ( .A(n277), .B(n278), .C(n279), .Z(n276) );
  GTECH_NOT U254 ( .A(n219), .Z(n221) );
  GTECH_NAND2 U255 ( .A(I_a[6]), .B(I_b[2]), .Z(n219) );
  GTECH_NOT U256 ( .A(n218), .Z(n222) );
  GTECH_NAND2 U257 ( .A(I_a[5]), .B(I_b[3]), .Z(n218) );
  GTECH_NOT U258 ( .A(n224), .Z(n267) );
  GTECH_OAI2N2 U259 ( .A(n280), .B(n281), .C(n282), .D(n283), .Z(n224) );
  GTECH_OR_NOT U260 ( .A(n284), .B(n280), .Z(n283) );
  GTECH_NOT U261 ( .A(n250), .Z(n251) );
  GTECH_OAI21 U262 ( .A(n285), .B(n286), .C(n287), .Z(n250) );
  GTECH_OAI21 U263 ( .A(n288), .B(n289), .C(n290), .Z(n287) );
  GTECH_XOR3 U264 ( .A(n291), .B(n286), .C(n289), .Z(N147) );
  GTECH_NOT U265 ( .A(n285), .Z(n289) );
  GTECH_XOR3 U266 ( .A(n292), .B(n281), .C(n280), .Z(n285) );
  GTECH_XOR3 U267 ( .A(n293), .B(n294), .C(n273), .Z(n280) );
  GTECH_OAI21 U268 ( .A(n295), .B(n296), .C(n297), .Z(n273) );
  GTECH_OAI21 U269 ( .A(n298), .B(n299), .C(n300), .Z(n297) );
  GTECH_NOT U270 ( .A(n271), .Z(n294) );
  GTECH_NAND2 U271 ( .A(I_a[7]), .B(I_b[0]), .Z(n271) );
  GTECH_NOT U272 ( .A(n270), .Z(n293) );
  GTECH_NAND2 U273 ( .A(I_a[6]), .B(I_b[1]), .Z(n270) );
  GTECH_NOT U274 ( .A(n284), .Z(n281) );
  GTECH_XOR3 U275 ( .A(n278), .B(n277), .C(n279), .Z(n284) );
  GTECH_OAI21 U276 ( .A(n301), .B(n302), .C(n303), .Z(n279) );
  GTECH_OAI21 U277 ( .A(n304), .B(n305), .C(n306), .Z(n303) );
  GTECH_NOT U278 ( .A(n275), .Z(n277) );
  GTECH_NAND2 U279 ( .A(I_a[5]), .B(I_b[2]), .Z(n275) );
  GTECH_NOT U280 ( .A(n274), .Z(n278) );
  GTECH_NAND2 U281 ( .A(I_a[4]), .B(I_b[3]), .Z(n274) );
  GTECH_NOT U282 ( .A(n282), .Z(n292) );
  GTECH_OAI2N2 U283 ( .A(n307), .B(n308), .C(n309), .D(n310), .Z(n282) );
  GTECH_OR_NOT U284 ( .A(n311), .B(n307), .Z(n310) );
  GTECH_NOT U285 ( .A(n288), .Z(n286) );
  GTECH_XOR3 U286 ( .A(n312), .B(n265), .C(n264), .Z(n288) );
  GTECH_XNOR2 U287 ( .A(n255), .B(n313), .Z(n264) );
  GTECH_AND2 U288 ( .A(I_b[7]), .B(I_a[0]), .Z(n313) );
  GTECH_NOT U289 ( .A(n314), .Z(n255) );
  GTECH_NAND2 U290 ( .A(I_b[6]), .B(I_a[1]), .Z(n314) );
  GTECH_NOT U291 ( .A(n266), .Z(n265) );
  GTECH_XOR3 U292 ( .A(n260), .B(n259), .C(n261), .Z(n266) );
  GTECH_OAI21 U293 ( .A(n315), .B(n316), .C(n317), .Z(n261) );
  GTECH_NOT U294 ( .A(n257), .Z(n259) );
  GTECH_NAND2 U295 ( .A(I_b[4]), .B(I_a[3]), .Z(n257) );
  GTECH_NOT U296 ( .A(n256), .Z(n260) );
  GTECH_NAND2 U297 ( .A(I_b[5]), .B(I_a[2]), .Z(n256) );
  GTECH_NOT U298 ( .A(n263), .Z(n312) );
  GTECH_NAND3 U299 ( .A(I_a[0]), .B(n318), .C(I_b[6]), .Z(n263) );
  GTECH_NOT U300 ( .A(n290), .Z(n291) );
  GTECH_OAI2N2 U301 ( .A(n319), .B(n320), .C(n321), .D(n322), .Z(n290) );
  GTECH_NAND2 U302 ( .A(n319), .B(n320), .Z(n322) );
  GTECH_XOR3 U303 ( .A(n323), .B(n324), .C(n319), .Z(N146) );
  GTECH_XOR3 U304 ( .A(n325), .B(n308), .C(n307), .Z(n319) );
  GTECH_XOR3 U305 ( .A(n295), .B(n296), .C(n300), .Z(n307) );
  GTECH_OAI21 U306 ( .A(n326), .B(n327), .C(n328), .Z(n300) );
  GTECH_OAI21 U307 ( .A(n329), .B(n330), .C(n331), .Z(n328) );
  GTECH_NOT U308 ( .A(n299), .Z(n296) );
  GTECH_NAND2 U309 ( .A(I_a[6]), .B(I_b[0]), .Z(n299) );
  GTECH_NOT U310 ( .A(n298), .Z(n295) );
  GTECH_NAND2 U311 ( .A(I_a[5]), .B(I_b[1]), .Z(n298) );
  GTECH_NOT U312 ( .A(n311), .Z(n308) );
  GTECH_XOR3 U313 ( .A(n305), .B(n304), .C(n306), .Z(n311) );
  GTECH_OAI21 U314 ( .A(n332), .B(n333), .C(n334), .Z(n306) );
  GTECH_OAI21 U315 ( .A(n335), .B(n336), .C(n337), .Z(n334) );
  GTECH_NOT U316 ( .A(n302), .Z(n304) );
  GTECH_NAND2 U317 ( .A(I_a[4]), .B(I_b[2]), .Z(n302) );
  GTECH_NOT U318 ( .A(n301), .Z(n305) );
  GTECH_NAND2 U319 ( .A(I_a[3]), .B(I_b[3]), .Z(n301) );
  GTECH_NOT U320 ( .A(n309), .Z(n325) );
  GTECH_OAI2N2 U321 ( .A(n338), .B(n339), .C(n340), .D(n341), .Z(n309) );
  GTECH_OR_NOT U322 ( .A(n342), .B(n338), .Z(n341) );
  GTECH_NOT U323 ( .A(n320), .Z(n324) );
  GTECH_XNOR2 U324 ( .A(n343), .B(n318), .Z(n320) );
  GTECH_NOT U325 ( .A(n344), .Z(n318) );
  GTECH_XOR3 U326 ( .A(n345), .B(n346), .C(n317), .Z(n344) );
  GTECH_NAND3 U327 ( .A(I_b[5]), .B(I_a[0]), .C(n347), .Z(n317) );
  GTECH_NOT U328 ( .A(n316), .Z(n346) );
  GTECH_NAND2 U329 ( .A(I_b[4]), .B(I_a[2]), .Z(n316) );
  GTECH_NOT U330 ( .A(n315), .Z(n345) );
  GTECH_NAND2 U331 ( .A(I_b[5]), .B(I_a[1]), .Z(n315) );
  GTECH_AND2 U332 ( .A(I_b[6]), .B(I_a[0]), .Z(n343) );
  GTECH_NOT U333 ( .A(n321), .Z(n323) );
  GTECH_OAI21 U334 ( .A(n348), .B(n349), .C(n350), .Z(n321) );
  GTECH_OAI21 U335 ( .A(n351), .B(n352), .C(n353), .Z(n350) );
  GTECH_XOR3 U336 ( .A(n353), .B(n351), .C(n352), .Z(N145) );
  GTECH_NOT U337 ( .A(n348), .Z(n352) );
  GTECH_XOR3 U338 ( .A(n354), .B(n339), .C(n338), .Z(n348) );
  GTECH_XOR3 U339 ( .A(n326), .B(n327), .C(n331), .Z(n338) );
  GTECH_OAI21 U340 ( .A(n355), .B(n356), .C(n357), .Z(n331) );
  GTECH_OAI21 U341 ( .A(n358), .B(n359), .C(n360), .Z(n357) );
  GTECH_NOT U342 ( .A(n330), .Z(n327) );
  GTECH_NAND2 U343 ( .A(I_a[5]), .B(I_b[0]), .Z(n330) );
  GTECH_NOT U344 ( .A(n329), .Z(n326) );
  GTECH_NAND2 U345 ( .A(I_a[4]), .B(I_b[1]), .Z(n329) );
  GTECH_NOT U346 ( .A(n342), .Z(n339) );
  GTECH_XOR3 U347 ( .A(n336), .B(n335), .C(n337), .Z(n342) );
  GTECH_OAI21 U348 ( .A(n361), .B(n362), .C(n363), .Z(n337) );
  GTECH_NOT U349 ( .A(n333), .Z(n335) );
  GTECH_NAND2 U350 ( .A(I_a[3]), .B(I_b[2]), .Z(n333) );
  GTECH_NOT U351 ( .A(n332), .Z(n336) );
  GTECH_NAND2 U352 ( .A(I_a[2]), .B(I_b[3]), .Z(n332) );
  GTECH_NOT U353 ( .A(n340), .Z(n354) );
  GTECH_OAI2N2 U354 ( .A(n364), .B(n365), .C(n366), .D(n367), .Z(n340) );
  GTECH_NAND2 U355 ( .A(n364), .B(n365), .Z(n367) );
  GTECH_NOT U356 ( .A(n349), .Z(n351) );
  GTECH_XNOR2 U357 ( .A(n347), .B(n368), .Z(n349) );
  GTECH_AND2 U358 ( .A(I_b[5]), .B(I_a[0]), .Z(n368) );
  GTECH_NOT U359 ( .A(n369), .Z(n347) );
  GTECH_NAND2 U360 ( .A(I_b[4]), .B(I_a[1]), .Z(n369) );
  GTECH_NOT U361 ( .A(n370), .Z(n353) );
  GTECH_NAND3 U362 ( .A(n371), .B(I_a[0]), .C(I_b[4]), .Z(n370) );
  GTECH_XNOR2 U363 ( .A(n371), .B(n372), .Z(N144) );
  GTECH_NAND2 U364 ( .A(I_b[4]), .B(I_a[0]), .Z(n372) );
  GTECH_XOR3 U365 ( .A(n373), .B(n374), .C(n364), .Z(n371) );
  GTECH_XOR3 U366 ( .A(n375), .B(n376), .C(n363), .Z(n364) );
  GTECH_NAND3 U367 ( .A(I_a[0]), .B(n377), .C(I_b[3]), .Z(n363) );
  GTECH_NOT U368 ( .A(n362), .Z(n376) );
  GTECH_NAND2 U369 ( .A(I_a[2]), .B(I_b[2]), .Z(n362) );
  GTECH_NOT U370 ( .A(n361), .Z(n375) );
  GTECH_NAND2 U371 ( .A(I_b[3]), .B(I_a[1]), .Z(n361) );
  GTECH_NOT U372 ( .A(n365), .Z(n374) );
  GTECH_XOR3 U373 ( .A(n355), .B(n356), .C(n360), .Z(n365) );
  GTECH_OAI22 U374 ( .A(n378), .B(n379), .C(n380), .D(n381), .Z(n360) );
  GTECH_NOR2 U375 ( .A(n382), .B(n383), .Z(n378) );
  GTECH_NOT U376 ( .A(n359), .Z(n356) );
  GTECH_NAND2 U377 ( .A(I_a[4]), .B(I_b[0]), .Z(n359) );
  GTECH_NOT U378 ( .A(n358), .Z(n355) );
  GTECH_NAND2 U379 ( .A(I_a[3]), .B(I_b[1]), .Z(n358) );
  GTECH_NOT U380 ( .A(n366), .Z(n373) );
  GTECH_OAI21 U381 ( .A(n384), .B(n385), .C(n386), .Z(n366) );
  GTECH_OAI21 U382 ( .A(n387), .B(n388), .C(n389), .Z(n386) );
  GTECH_NOT U383 ( .A(n388), .Z(n384) );
  GTECH_XOR3 U384 ( .A(n389), .B(n387), .C(n388), .Z(N143) );
  GTECH_XOR3 U385 ( .A(n380), .B(n381), .C(n379), .Z(n388) );
  GTECH_OAI21 U386 ( .A(n390), .B(n391), .C(n392), .Z(n379) );
  GTECH_NOT U387 ( .A(n383), .Z(n381) );
  GTECH_NAND2 U388 ( .A(I_a[3]), .B(I_b[0]), .Z(n383) );
  GTECH_NOT U389 ( .A(n382), .Z(n380) );
  GTECH_NAND2 U390 ( .A(I_b[1]), .B(I_a[2]), .Z(n382) );
  GTECH_NOT U391 ( .A(n385), .Z(n387) );
  GTECH_XNOR2 U392 ( .A(n377), .B(n393), .Z(n385) );
  GTECH_AND2 U393 ( .A(I_b[3]), .B(I_a[0]), .Z(n393) );
  GTECH_NOT U394 ( .A(n394), .Z(n377) );
  GTECH_NAND2 U395 ( .A(I_b[2]), .B(I_a[1]), .Z(n394) );
  GTECH_NOT U396 ( .A(n395), .Z(n389) );
  GTECH_NAND3 U397 ( .A(I_b[2]), .B(n396), .C(I_a[0]), .Z(n395) );
  GTECH_NOT U398 ( .A(n397), .Z(n396) );
  GTECH_XNOR2 U399 ( .A(n398), .B(n397), .Z(N142) );
  GTECH_XOR3 U400 ( .A(n399), .B(n400), .C(n392), .Z(n397) );
  GTECH_NAND3 U401 ( .A(n401), .B(I_a[0]), .C(I_b[1]), .Z(n392) );
  GTECH_NOT U402 ( .A(n391), .Z(n400) );
  GTECH_NAND2 U403 ( .A(I_b[0]), .B(I_a[2]), .Z(n391) );
  GTECH_NOT U404 ( .A(n390), .Z(n399) );
  GTECH_NAND2 U405 ( .A(I_b[1]), .B(I_a[1]), .Z(n390) );
  GTECH_AND2 U406 ( .A(I_a[0]), .B(I_b[2]), .Z(n398) );
  GTECH_XNOR2 U407 ( .A(n401), .B(n402), .Z(N141) );
  GTECH_NAND2 U408 ( .A(I_b[1]), .B(I_a[0]), .Z(n402) );
  GTECH_NOT U409 ( .A(n403), .Z(n401) );
  GTECH_NAND2 U410 ( .A(I_b[0]), .B(I_a[1]), .Z(n403) );
  GTECH_AND2 U411 ( .A(I_b[0]), .B(I_a[0]), .Z(N140) );
endmodule

