
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379;

  GTECH_MUX2 U134 ( .A(n273), .B(n274), .S(n275), .Z(sum[9]) );
  GTECH_AOI21 U135 ( .A(n276), .B(n277), .C(n278), .Z(n275) );
  GTECH_XOR2 U136 ( .A(b[9]), .B(a[9]), .Z(n274) );
  GTECH_OR_NOT U137 ( .A(n279), .B(n280), .Z(n273) );
  GTECH_XNOR2 U138 ( .A(n281), .B(n282), .Z(sum[8]) );
  GTECH_MUX2 U139 ( .A(n283), .B(n284), .S(n285), .Z(sum[7]) );
  GTECH_XNOR2 U140 ( .A(n286), .B(n287), .Z(n284) );
  GTECH_AND_NOT U141 ( .A(n288), .B(n289), .Z(n287) );
  GTECH_OAI21 U142 ( .A(b[6]), .B(a[6]), .C(n290), .Z(n288) );
  GTECH_XOR2 U143 ( .A(n286), .B(n291), .Z(n283) );
  GTECH_XOR2 U144 ( .A(a[7]), .B(b[7]), .Z(n286) );
  GTECH_AO21 U145 ( .A(n292), .B(n289), .C(n293), .Z(sum[6]) );
  GTECH_NOT U146 ( .A(n294), .Z(n293) );
  GTECH_MUX2 U147 ( .A(n295), .B(n296), .S(b[6]), .Z(n294) );
  GTECH_OR2 U148 ( .A(n292), .B(a[6]), .Z(n296) );
  GTECH_XNOR2 U149 ( .A(a[6]), .B(n292), .Z(n295) );
  GTECH_AO21 U150 ( .A(n297), .B(n298), .C(n290), .Z(n292) );
  GTECH_OAI21 U151 ( .A(n299), .B(n300), .C(n301), .Z(n290) );
  GTECH_MUX2 U152 ( .A(n302), .B(n303), .S(n304), .Z(sum[5]) );
  GTECH_AND_NOT U153 ( .A(n301), .B(n299), .Z(n304) );
  GTECH_OAI21 U154 ( .A(a[4]), .B(n298), .C(n305), .Z(n303) );
  GTECH_AO21 U155 ( .A(n298), .B(a[4]), .C(b[4]), .Z(n305) );
  GTECH_OAI21 U156 ( .A(n306), .B(n285), .C(n300), .Z(n302) );
  GTECH_XNOR2 U157 ( .A(n285), .B(n307), .Z(sum[4]) );
  GTECH_MUX2 U158 ( .A(n308), .B(n309), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U159 ( .A(n310), .B(n311), .Z(n309) );
  GTECH_XOR2 U160 ( .A(n312), .B(n310), .Z(n308) );
  GTECH_XOR2 U161 ( .A(a[3]), .B(b[3]), .Z(n310) );
  GTECH_OA21 U162 ( .A(a[2]), .B(n313), .C(n314), .Z(n312) );
  GTECH_AO21 U163 ( .A(n313), .B(a[2]), .C(b[2]), .Z(n314) );
  GTECH_MUX2 U164 ( .A(n315), .B(n316), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U165 ( .A(n317), .B(n318), .Z(n316) );
  GTECH_XNOR2 U166 ( .A(n317), .B(n313), .Z(n315) );
  GTECH_OAI21 U167 ( .A(n319), .B(n320), .C(n321), .Z(n313) );
  GTECH_XNOR2 U168 ( .A(a[2]), .B(b[2]), .Z(n317) );
  GTECH_MUX2 U169 ( .A(n322), .B(n323), .S(n324), .Z(sum[1]) );
  GTECH_AND_NOT U170 ( .A(n321), .B(n319), .Z(n324) );
  GTECH_AO21 U171 ( .A(n325), .B(n320), .C(n326), .Z(n323) );
  GTECH_OAI21 U172 ( .A(n326), .B(n325), .C(n320), .Z(n322) );
  GTECH_OR_NOT U173 ( .A(n327), .B(b[0]), .Z(n320) );
  GTECH_NOT U174 ( .A(cin), .Z(n325) );
  GTECH_MUX2 U175 ( .A(n328), .B(n329), .S(n330), .Z(sum[15]) );
  GTECH_XNOR2 U176 ( .A(n331), .B(n332), .Z(n329) );
  GTECH_XOR2 U177 ( .A(n331), .B(n333), .Z(n328) );
  GTECH_AND_NOT U178 ( .A(n334), .B(n335), .Z(n333) );
  GTECH_OAI21 U179 ( .A(b[14]), .B(a[14]), .C(n336), .Z(n334) );
  GTECH_XNOR2 U180 ( .A(a[15]), .B(b[15]), .Z(n331) );
  GTECH_AO21 U181 ( .A(n337), .B(n335), .C(n338), .Z(sum[14]) );
  GTECH_NOT U182 ( .A(n339), .Z(n338) );
  GTECH_MUX2 U183 ( .A(n340), .B(n341), .S(b[14]), .Z(n339) );
  GTECH_OR2 U184 ( .A(a[14]), .B(n337), .Z(n341) );
  GTECH_XNOR2 U185 ( .A(a[14]), .B(n337), .Z(n340) );
  GTECH_AO21 U186 ( .A(n342), .B(n330), .C(n336), .Z(n337) );
  GTECH_AO22 U187 ( .A(a[13]), .B(b[13]), .C(n343), .D(n344), .Z(n336) );
  GTECH_MUX2 U188 ( .A(n345), .B(n346), .S(n330), .Z(sum[13]) );
  GTECH_XOR2 U189 ( .A(n347), .B(n348), .Z(n346) );
  GTECH_XOR2 U190 ( .A(n348), .B(n344), .Z(n345) );
  GTECH_AOI21 U191 ( .A(a[13]), .B(b[13]), .C(n349), .Z(n348) );
  GTECH_NOT U192 ( .A(n343), .Z(n349) );
  GTECH_XNOR2 U193 ( .A(n350), .B(n330), .Z(sum[12]) );
  GTECH_MUX2 U194 ( .A(n351), .B(n352), .S(n281), .Z(sum[11]) );
  GTECH_XNOR2 U195 ( .A(n353), .B(n354), .Z(n352) );
  GTECH_OA21 U196 ( .A(a[10]), .B(n355), .C(n356), .Z(n353) );
  GTECH_AO21 U197 ( .A(n355), .B(a[10]), .C(b[10]), .Z(n356) );
  GTECH_XNOR2 U198 ( .A(n354), .B(n357), .Z(n351) );
  GTECH_XNOR2 U199 ( .A(a[11]), .B(b[11]), .Z(n354) );
  GTECH_MUX2 U200 ( .A(n358), .B(n359), .S(n281), .Z(sum[10]) );
  GTECH_NOT U201 ( .A(n277), .Z(n281) );
  GTECH_XNOR2 U202 ( .A(n360), .B(n355), .Z(n359) );
  GTECH_AO21 U203 ( .A(n280), .B(n278), .C(n279), .Z(n355) );
  GTECH_XNOR2 U204 ( .A(n360), .B(n361), .Z(n358) );
  GTECH_XNOR2 U205 ( .A(a[10]), .B(b[10]), .Z(n360) );
  GTECH_XOR2 U206 ( .A(cin), .B(n362), .Z(sum[0]) );
  GTECH_NOT U207 ( .A(n363), .Z(cout) );
  GTECH_MUX2 U208 ( .A(n350), .B(n364), .S(n330), .Z(n363) );
  GTECH_MUX2 U209 ( .A(n282), .B(n365), .S(n277), .Z(n330) );
  GTECH_MUX2 U210 ( .A(n366), .B(n307), .S(n285), .Z(n277) );
  GTECH_NOT U211 ( .A(n298), .Z(n285) );
  GTECH_MUX2 U212 ( .A(n362), .B(n367), .S(cin), .Z(n298) );
  GTECH_OA21 U213 ( .A(a[3]), .B(n311), .C(n368), .Z(n367) );
  GTECH_AO21 U214 ( .A(n311), .B(a[3]), .C(b[3]), .Z(n368) );
  GTECH_AO21 U215 ( .A(n318), .B(a[2]), .C(n369), .Z(n311) );
  GTECH_OA21 U216 ( .A(a[2]), .B(n318), .C(b[2]), .Z(n369) );
  GTECH_OAI21 U217 ( .A(n326), .B(n319), .C(n321), .Z(n318) );
  GTECH_OR_NOT U218 ( .A(n370), .B(a[1]), .Z(n321) );
  GTECH_AND_NOT U219 ( .A(n370), .B(a[1]), .Z(n319) );
  GTECH_NOT U220 ( .A(b[1]), .Z(n370) );
  GTECH_AND2 U221 ( .A(n327), .B(n371), .Z(n326) );
  GTECH_XOR2 U222 ( .A(n327), .B(n371), .Z(n362) );
  GTECH_NOT U223 ( .A(b[0]), .Z(n371) );
  GTECH_NOT U224 ( .A(a[0]), .Z(n327) );
  GTECH_AND_NOT U225 ( .A(n300), .B(n306), .Z(n307) );
  GTECH_OR_NOT U226 ( .A(n372), .B(b[4]), .Z(n300) );
  GTECH_OA21 U227 ( .A(a[7]), .B(n291), .C(n373), .Z(n366) );
  GTECH_AO21 U228 ( .A(n291), .B(a[7]), .C(b[7]), .Z(n373) );
  GTECH_AO21 U229 ( .A(n297), .B(n374), .C(n289), .Z(n291) );
  GTECH_AND2 U230 ( .A(b[6]), .B(a[6]), .Z(n289) );
  GTECH_OR2 U231 ( .A(b[6]), .B(a[6]), .Z(n374) );
  GTECH_OAI21 U232 ( .A(n306), .B(n299), .C(n301), .Z(n297) );
  GTECH_OR_NOT U233 ( .A(n375), .B(b[5]), .Z(n301) );
  GTECH_AND_NOT U234 ( .A(n375), .B(b[5]), .Z(n299) );
  GTECH_NOT U235 ( .A(a[5]), .Z(n375) );
  GTECH_AND_NOT U236 ( .A(n372), .B(b[4]), .Z(n306) );
  GTECH_NOT U237 ( .A(a[4]), .Z(n372) );
  GTECH_AO21 U238 ( .A(n357), .B(a[11]), .C(n376), .Z(n365) );
  GTECH_OA21 U239 ( .A(a[11]), .B(n357), .C(b[11]), .Z(n376) );
  GTECH_AO21 U240 ( .A(n361), .B(a[10]), .C(n377), .Z(n357) );
  GTECH_OA21 U241 ( .A(a[10]), .B(n361), .C(b[10]), .Z(n377) );
  GTECH_AO21 U242 ( .A(n276), .B(n280), .C(n279), .Z(n361) );
  GTECH_AND2 U243 ( .A(a[9]), .B(b[9]), .Z(n279) );
  GTECH_OR2 U244 ( .A(a[9]), .B(b[9]), .Z(n280) );
  GTECH_AND_NOT U245 ( .A(n276), .B(n278), .Z(n282) );
  GTECH_AND2 U246 ( .A(b[8]), .B(a[8]), .Z(n278) );
  GTECH_OR2 U247 ( .A(a[8]), .B(b[8]), .Z(n276) );
  GTECH_AOI21 U248 ( .A(n332), .B(a[15]), .C(n378), .Z(n364) );
  GTECH_OA21 U249 ( .A(a[15]), .B(n332), .C(b[15]), .Z(n378) );
  GTECH_AO21 U250 ( .A(n342), .B(n379), .C(n335), .Z(n332) );
  GTECH_AND2 U251 ( .A(b[14]), .B(a[14]), .Z(n335) );
  GTECH_OR2 U252 ( .A(b[14]), .B(a[14]), .Z(n379) );
  GTECH_AO22 U253 ( .A(a[13]), .B(b[13]), .C(n347), .D(n343), .Z(n342) );
  GTECH_OR2 U254 ( .A(a[13]), .B(b[13]), .Z(n343) );
  GTECH_OR_NOT U255 ( .A(n344), .B(n347), .Z(n350) );
  GTECH_OR2 U256 ( .A(a[12]), .B(b[12]), .Z(n347) );
  GTECH_AND2 U257 ( .A(b[12]), .B(a[12]), .Z(n344) );
endmodule

