
module CRC32 ( crcIn, data, crcOut );
  input [31:0] crcIn;
  input [7:0] data;
  output [31:0] crcOut;
  wire   n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58;

  GTECH_XOR2 U62 ( .A(crcIn[17]), .B(n30), .Z(crcOut[9]) );
  GTECH_XOR3 U63 ( .A(crcIn[16]), .B(n31), .C(n32), .Z(crcOut[8]) );
  GTECH_XOR3 U64 ( .A(crcIn[15]), .B(n33), .C(n34), .Z(crcOut[7]) );
  GTECH_NOT U65 ( .A(n35), .Z(n33) );
  GTECH_XOR2 U66 ( .A(crcIn[14]), .B(n36), .Z(crcOut[6]) );
  GTECH_XNOR3 U67 ( .A(crcIn[13]), .B(crcOut[31]), .C(n37), .Z(crcOut[5]) );
  GTECH_XNOR3 U68 ( .A(crcIn[12]), .B(n35), .C(n38), .Z(crcOut[4]) );
  GTECH_XNOR3 U69 ( .A(crcIn[11]), .B(n39), .C(n40), .Z(crcOut[3]) );
  GTECH_XOR3 U70 ( .A(crcIn[10]), .B(n41), .C(n42), .Z(crcOut[2]) );
  GTECH_XOR2 U71 ( .A(n34), .B(crcOut[30]), .Z(crcOut[29]) );
  GTECH_XNOR2 U72 ( .A(n35), .B(n36), .Z(crcOut[28]) );
  GTECH_XOR2 U73 ( .A(n43), .B(n44), .Z(n35) );
  GTECH_XOR3 U74 ( .A(n36), .B(crcOut[31]), .C(n45), .Z(crcOut[27]) );
  GTECH_XNOR2 U75 ( .A(n31), .B(n46), .Z(crcOut[31]) );
  GTECH_XOR3 U76 ( .A(n41), .B(n38), .C(crcOut[30]), .Z(crcOut[26]) );
  GTECH_XOR2 U77 ( .A(n42), .B(n32), .Z(crcOut[30]) );
  GTECH_XOR2 U78 ( .A(n42), .B(n47), .Z(crcOut[25]) );
  GTECH_XOR2 U79 ( .A(n43), .B(n48), .Z(crcOut[24]) );
  GTECH_XNOR2 U80 ( .A(crcIn[31]), .B(n49), .Z(crcOut[23]) );
  GTECH_XOR2 U81 ( .A(crcIn[30]), .B(n47), .Z(crcOut[22]) );
  GTECH_XOR3 U82 ( .A(n44), .B(n50), .C(n38), .Z(n47) );
  GTECH_XOR2 U83 ( .A(crcIn[29]), .B(n48), .Z(crcOut[21]) );
  GTECH_XOR3 U84 ( .A(n30), .B(n36), .C(n39), .Z(n48) );
  GTECH_XNOR2 U85 ( .A(crcIn[28]), .B(n49), .Z(crcOut[20]) );
  GTECH_XOR2 U86 ( .A(n37), .B(n32), .Z(n49) );
  GTECH_XOR2 U87 ( .A(n45), .B(n51), .Z(n37) );
  GTECH_XOR3 U88 ( .A(crcIn[9]), .B(n43), .C(n45), .Z(crcOut[1]) );
  GTECH_XOR4 U89 ( .A(n52), .B(n40), .C(crcIn[27]), .D(n32), .Z(crcOut[19]) );
  GTECH_XOR2 U90 ( .A(n53), .B(n30), .Z(n32) );
  GTECH_NOT U91 ( .A(n46), .Z(n30) );
  GTECH_XOR2 U92 ( .A(n50), .B(n31), .Z(n40) );
  GTECH_XOR3 U93 ( .A(crcIn[26]), .B(n54), .C(n55), .Z(crcOut[18]) );
  GTECH_XNOR3 U94 ( .A(crcIn[25]), .B(n45), .C(n54), .Z(crcOut[17]) );
  GTECH_XNOR2 U95 ( .A(n42), .B(n36), .Z(n54) );
  GTECH_XNOR2 U96 ( .A(n41), .B(n50), .Z(n36) );
  GTECH_NOT U97 ( .A(n51), .Z(n41) );
  GTECH_XOR3 U98 ( .A(crcIn[24]), .B(n52), .C(n56), .Z(crcOut[16]) );
  GTECH_NOT U99 ( .A(n38), .Z(n52) );
  GTECH_XNOR3 U100 ( .A(crcIn[23]), .B(n46), .C(n38), .Z(crcOut[15]) );
  GTECH_XNOR2 U101 ( .A(n57), .B(n45), .Z(n38) );
  GTECH_XNOR2 U102 ( .A(data[7]), .B(crcIn[7]), .Z(n46) );
  GTECH_XNOR3 U103 ( .A(crcIn[22]), .B(n31), .C(n55), .Z(crcOut[14]) );
  GTECH_XOR2 U104 ( .A(n57), .B(n53), .Z(n55) );
  GTECH_NOT U105 ( .A(n44), .Z(n53) );
  GTECH_XNOR2 U106 ( .A(data[6]), .B(crcIn[6]), .Z(n44) );
  GTECH_NOT U107 ( .A(n58), .Z(n31) );
  GTECH_XOR3 U108 ( .A(crcIn[21]), .B(n34), .C(n42), .Z(crcOut[13]) );
  GTECH_XNOR2 U109 ( .A(n43), .B(n58), .Z(n42) );
  GTECH_XNOR2 U110 ( .A(data[1]), .B(crcIn[1]), .Z(n58) );
  GTECH_NOT U111 ( .A(n50), .Z(n34) );
  GTECH_XNOR2 U112 ( .A(data[5]), .B(crcIn[5]), .Z(n50) );
  GTECH_XNOR2 U113 ( .A(crcIn[20]), .B(n56), .Z(crcOut[12]) );
  GTECH_XOR2 U114 ( .A(n51), .B(n43), .Z(n56) );
  GTECH_XOR2 U115 ( .A(data[0]), .B(crcIn[0]), .Z(n43) );
  GTECH_XNOR2 U116 ( .A(data[4]), .B(crcIn[4]), .Z(n51) );
  GTECH_XOR2 U117 ( .A(crcIn[19]), .B(n45), .Z(crcOut[11]) );
  GTECH_XOR2 U118 ( .A(data[3]), .B(crcIn[3]), .Z(n45) );
  GTECH_XOR2 U119 ( .A(crcIn[18]), .B(n39), .Z(crcOut[10]) );
  GTECH_XOR2 U120 ( .A(crcIn[8]), .B(n39), .Z(crcOut[0]) );
  GTECH_NOT U121 ( .A(n57), .Z(n39) );
  GTECH_XNOR2 U122 ( .A(data[2]), .B(crcIn[2]), .Z(n57) );
endmodule

