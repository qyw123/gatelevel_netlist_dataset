
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375;

  GTECH_OAI22 U132 ( .A(n271), .B(n272), .C(n273), .D(n274), .Z(sum[9]) );
  GTECH_XNOR2 U133 ( .A(n275), .B(n276), .Z(n274) );
  GTECH_XOR2 U134 ( .A(n275), .B(n277), .Z(n271) );
  GTECH_AOI21 U135 ( .A(n278), .B(n279), .C(n280), .Z(n275) );
  GTECH_OR_NOT U136 ( .A(n281), .B(n282), .Z(sum[8]) );
  GTECH_OAI21 U137 ( .A(n276), .B(n277), .C(n273), .Z(n282) );
  GTECH_OAI22 U138 ( .A(n283), .B(n284), .C(n285), .D(n286), .Z(sum[7]) );
  GTECH_XNOR2 U139 ( .A(n287), .B(n288), .Z(n286) );
  GTECH_AOI2N2 U140 ( .A(n289), .B(n290), .C(b[6]), .D(n291), .Z(n288) );
  GTECH_NOR2 U141 ( .A(n289), .B(n290), .Z(n291) );
  GTECH_XNOR2 U142 ( .A(n292), .B(n287), .Z(n283) );
  GTECH_XOR2 U143 ( .A(a[7]), .B(b[7]), .Z(n287) );
  GTECH_OAI22 U144 ( .A(n293), .B(n284), .C(n294), .D(n285), .Z(sum[6]) );
  GTECH_XOR2 U145 ( .A(n290), .B(n295), .Z(n294) );
  GTECH_AOI21 U146 ( .A(n296), .B(n297), .C(n298), .Z(n290) );
  GTECH_XNOR2 U147 ( .A(n299), .B(n295), .Z(n293) );
  GTECH_XNOR2 U148 ( .A(n289), .B(b[6]), .Z(n295) );
  GTECH_NOT U149 ( .A(a[6]), .Z(n289) );
  GTECH_OAI2N2 U150 ( .A(n300), .B(n301), .C(n302), .D(n300), .Z(sum[5]) );
  GTECH_OAI21 U151 ( .A(n285), .B(n297), .C(n303), .Z(n302) );
  GTECH_AOI21 U152 ( .A(n285), .B(n303), .C(n297), .Z(n301) );
  GTECH_AND2 U153 ( .A(a[4]), .B(b[4]), .Z(n297) );
  GTECH_AND_NOT U154 ( .A(n296), .B(n298), .Z(n300) );
  GTECH_XNOR2 U155 ( .A(n284), .B(n304), .Z(sum[4]) );
  GTECH_OAI22 U156 ( .A(n305), .B(n306), .C(cin), .D(n307), .Z(sum[3]) );
  GTECH_XNOR2 U157 ( .A(n308), .B(n309), .Z(n307) );
  GTECH_AOI21 U158 ( .A(n310), .B(n311), .C(n312), .Z(n309) );
  GTECH_XNOR2 U159 ( .A(n308), .B(n313), .Z(n306) );
  GTECH_XOR2 U160 ( .A(a[3]), .B(b[3]), .Z(n308) );
  GTECH_OAI22 U161 ( .A(n305), .B(n314), .C(cin), .D(n315), .Z(sum[2]) );
  GTECH_XNOR2 U162 ( .A(n316), .B(n310), .Z(n315) );
  GTECH_AOI21 U163 ( .A(n317), .B(n318), .C(n319), .Z(n310) );
  GTECH_XNOR2 U164 ( .A(n320), .B(n316), .Z(n314) );
  GTECH_OAI21 U165 ( .A(a[2]), .B(b[2]), .C(n311), .Z(n316) );
  GTECH_OAI2N2 U166 ( .A(n321), .B(n322), .C(n323), .D(n322), .Z(sum[1]) );
  GTECH_AO21 U167 ( .A(cin), .B(n324), .C(n318), .Z(n323) );
  GTECH_NOT U168 ( .A(n325), .Z(n318) );
  GTECH_OR_NOT U169 ( .A(n319), .B(n317), .Z(n322) );
  GTECH_AOI21 U170 ( .A(n325), .B(n305), .C(n326), .Z(n321) );
  GTECH_OAI22 U171 ( .A(n327), .B(n328), .C(n329), .D(n330), .Z(sum[15]) );
  GTECH_XNOR2 U172 ( .A(n331), .B(n332), .Z(n330) );
  GTECH_XNOR2 U173 ( .A(n333), .B(n332), .Z(n328) );
  GTECH_XOR2 U174 ( .A(a[15]), .B(b[15]), .Z(n332) );
  GTECH_OAI21 U175 ( .A(n334), .B(n335), .C(n336), .Z(n333) );
  GTECH_OAI22 U176 ( .A(n327), .B(n337), .C(n329), .D(n338), .Z(sum[14]) );
  GTECH_XOR2 U177 ( .A(n339), .B(n340), .Z(n338) );
  GTECH_XOR2 U178 ( .A(n340), .B(n334), .Z(n337) );
  GTECH_AOI21 U179 ( .A(n341), .B(n342), .C(n343), .Z(n334) );
  GTECH_AND_NOT U180 ( .A(n336), .B(n335), .Z(n340) );
  GTECH_OAI22 U181 ( .A(n327), .B(n344), .C(n329), .D(n345), .Z(sum[13]) );
  GTECH_XOR2 U182 ( .A(n346), .B(n347), .Z(n345) );
  GTECH_NOT U183 ( .A(n327), .Z(n329) );
  GTECH_XOR2 U184 ( .A(n347), .B(n342), .Z(n344) );
  GTECH_OR_NOT U185 ( .A(n343), .B(n341), .Z(n347) );
  GTECH_OR_NOT U186 ( .A(n348), .B(n349), .Z(sum[12]) );
  GTECH_OAI21 U187 ( .A(n342), .B(n350), .C(n327), .Z(n349) );
  GTECH_OAI22 U188 ( .A(n273), .B(n351), .C(n272), .D(n352), .Z(sum[11]) );
  GTECH_XNOR2 U189 ( .A(n353), .B(n354), .Z(n352) );
  GTECH_XOR2 U190 ( .A(n353), .B(n355), .Z(n351) );
  GTECH_AO21 U191 ( .A(n356), .B(n357), .C(n358), .Z(n355) );
  GTECH_XOR2 U192 ( .A(a[11]), .B(b[11]), .Z(n353) );
  GTECH_OAI22 U193 ( .A(n359), .B(n272), .C(n360), .D(n273), .Z(sum[10]) );
  GTECH_XNOR2 U194 ( .A(n361), .B(n356), .Z(n360) );
  GTECH_AND_NOT U195 ( .A(n362), .B(n280), .Z(n356) );
  GTECH_OAI21 U196 ( .A(a[9]), .B(b[9]), .C(n276), .Z(n362) );
  GTECH_XNOR2 U197 ( .A(n363), .B(n361), .Z(n359) );
  GTECH_OAI21 U198 ( .A(a[10]), .B(b[10]), .C(n357), .Z(n361) );
  GTECH_XOR2 U199 ( .A(n305), .B(n364), .Z(sum[0]) );
  GTECH_AO21 U200 ( .A(n327), .B(n365), .C(n348), .Z(cout) );
  GTECH_NOR3 U201 ( .A(n342), .B(n350), .C(n327), .Z(n348) );
  GTECH_NOT U202 ( .A(n346), .Z(n350) );
  GTECH_AND2 U203 ( .A(b[12]), .B(a[12]), .Z(n342) );
  GTECH_AO22 U204 ( .A(n366), .B(b[15]), .C(n331), .D(a[15]), .Z(n365) );
  GTECH_NOT U205 ( .A(n367), .Z(n366) );
  GTECH_NOR2 U206 ( .A(n331), .B(a[15]), .Z(n367) );
  GTECH_OAI21 U207 ( .A(n339), .B(n335), .C(n336), .Z(n331) );
  GTECH_NAND2 U208 ( .A(a[14]), .B(b[14]), .Z(n336) );
  GTECH_NOR2 U209 ( .A(b[14]), .B(a[14]), .Z(n335) );
  GTECH_AOI21 U210 ( .A(n341), .B(n346), .C(n343), .Z(n339) );
  GTECH_AND2 U211 ( .A(b[13]), .B(a[13]), .Z(n343) );
  GTECH_OR2 U212 ( .A(a[12]), .B(b[12]), .Z(n346) );
  GTECH_OR2 U213 ( .A(a[13]), .B(b[13]), .Z(n341) );
  GTECH_AO21 U214 ( .A(n273), .B(n368), .C(n281), .Z(n327) );
  GTECH_NOR3 U215 ( .A(n277), .B(n276), .C(n273), .Z(n281) );
  GTECH_AND2 U216 ( .A(a[8]), .B(b[8]), .Z(n276) );
  GTECH_ADD_ABC U217 ( .A(n354), .B(a[11]), .C(b[11]), .COUT(n368) );
  GTECH_AOI21 U218 ( .A(n357), .B(n363), .C(n358), .Z(n354) );
  GTECH_NOR2 U219 ( .A(b[10]), .B(a[10]), .Z(n358) );
  GTECH_AND_NOT U220 ( .A(n369), .B(n280), .Z(n363) );
  GTECH_AND_NOT U221 ( .A(a[9]), .B(n278), .Z(n280) );
  GTECH_AO21 U222 ( .A(n278), .B(n279), .C(n277), .Z(n369) );
  GTECH_NOR2 U223 ( .A(b[8]), .B(a[8]), .Z(n277) );
  GTECH_NOT U224 ( .A(a[9]), .Z(n279) );
  GTECH_NOT U225 ( .A(b[9]), .Z(n278) );
  GTECH_NAND2 U226 ( .A(a[10]), .B(b[10]), .Z(n357) );
  GTECH_NOT U227 ( .A(n272), .Z(n273) );
  GTECH_OAI22 U228 ( .A(n370), .B(n284), .C(n304), .D(n285), .Z(n272) );
  GTECH_NOT U229 ( .A(n284), .Z(n285) );
  GTECH_XNOR2 U230 ( .A(a[4]), .B(n371), .Z(n304) );
  GTECH_NOT U231 ( .A(b[4]), .Z(n371) );
  GTECH_OAI2N2 U232 ( .A(n372), .B(n305), .C(n305), .D(n364), .Z(n284) );
  GTECH_NAND2 U233 ( .A(n324), .B(n325), .Z(n364) );
  GTECH_NAND2 U234 ( .A(b[0]), .B(a[0]), .Z(n325) );
  GTECH_NOT U235 ( .A(cin), .Z(n305) );
  GTECH_ADD_ABC U236 ( .A(a[3]), .B(n313), .C(b[3]), .COUT(n372) );
  GTECH_AOI21 U237 ( .A(n311), .B(n320), .C(n312), .Z(n313) );
  GTECH_NOR2 U238 ( .A(b[2]), .B(a[2]), .Z(n312) );
  GTECH_AOI21 U239 ( .A(n324), .B(n317), .C(n319), .Z(n320) );
  GTECH_AND2 U240 ( .A(b[1]), .B(a[1]), .Z(n319) );
  GTECH_OR2 U241 ( .A(a[1]), .B(b[1]), .Z(n317) );
  GTECH_NOT U242 ( .A(n326), .Z(n324) );
  GTECH_NOR2 U243 ( .A(a[0]), .B(b[0]), .Z(n326) );
  GTECH_NAND2 U244 ( .A(a[2]), .B(b[2]), .Z(n311) );
  GTECH_OA22 U245 ( .A(b[7]), .B(n373), .C(a[7]), .D(n292), .Z(n370) );
  GTECH_AND2 U246 ( .A(n292), .B(a[7]), .Z(n373) );
  GTECH_AO21 U247 ( .A(n299), .B(a[6]), .C(n374), .Z(n292) );
  GTECH_NOT U248 ( .A(n375), .Z(n374) );
  GTECH_OAI21 U249 ( .A(a[6]), .B(n299), .C(b[6]), .Z(n375) );
  GTECH_AO21 U250 ( .A(n303), .B(n296), .C(n298), .Z(n299) );
  GTECH_AND2 U251 ( .A(b[5]), .B(a[5]), .Z(n298) );
  GTECH_OR2 U252 ( .A(a[5]), .B(b[5]), .Z(n296) );
  GTECH_OR2 U253 ( .A(a[4]), .B(b[4]), .Z(n303) );
endmodule

