
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387;

  GTECH_MUX2 U139 ( .A(n278), .B(n279), .S(n280), .Z(sum[9]) );
  GTECH_AOI21 U140 ( .A(n281), .B(n282), .C(n283), .Z(n280) );
  GTECH_OR_NOT U141 ( .A(n284), .B(n285), .Z(n279) );
  GTECH_XOR2 U142 ( .A(b[9]), .B(a[9]), .Z(n278) );
  GTECH_NAND2 U143 ( .A(n286), .B(n287), .Z(sum[8]) );
  GTECH_AO21 U144 ( .A(n288), .B(n281), .C(n282), .Z(n286) );
  GTECH_MUX2 U145 ( .A(n289), .B(n290), .S(n291), .Z(sum[7]) );
  GTECH_XOR2 U146 ( .A(n292), .B(n293), .Z(n290) );
  GTECH_XNOR2 U147 ( .A(n292), .B(n294), .Z(n289) );
  GTECH_OA21 U148 ( .A(n295), .B(n296), .C(n297), .Z(n294) );
  GTECH_NOR2 U149 ( .A(b[6]), .B(a[6]), .Z(n295) );
  GTECH_XOR2 U150 ( .A(a[7]), .B(b[7]), .Z(n292) );
  GTECH_OAI21 U151 ( .A(n298), .B(n297), .C(n299), .Z(sum[6]) );
  GTECH_MUX2 U152 ( .A(n300), .B(n301), .S(b[6]), .Z(n299) );
  GTECH_OR_NOT U153 ( .A(a[6]), .B(n298), .Z(n301) );
  GTECH_XOR2 U154 ( .A(a[6]), .B(n298), .Z(n300) );
  GTECH_AOI21 U155 ( .A(n291), .B(n302), .C(n303), .Z(n298) );
  GTECH_NOT U156 ( .A(n296), .Z(n303) );
  GTECH_OAI21 U157 ( .A(n304), .B(n305), .C(n306), .Z(n296) );
  GTECH_MUX2 U158 ( .A(n307), .B(n308), .S(n309), .Z(sum[5]) );
  GTECH_AND_NOT U159 ( .A(n306), .B(n305), .Z(n309) );
  GTECH_OAI21 U160 ( .A(n304), .B(n291), .C(n310), .Z(n308) );
  GTECH_AO21 U161 ( .A(n310), .B(n291), .C(n304), .Z(n307) );
  GTECH_XNOR2 U162 ( .A(n311), .B(n312), .Z(sum[4]) );
  GTECH_MUX2 U163 ( .A(n313), .B(n314), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U164 ( .A(n315), .B(n316), .Z(n314) );
  GTECH_XNOR2 U165 ( .A(n315), .B(n317), .Z(n313) );
  GTECH_OA21 U166 ( .A(n318), .B(n319), .C(n320), .Z(n317) );
  GTECH_NOR2 U167 ( .A(a[2]), .B(b[2]), .Z(n318) );
  GTECH_XOR2 U168 ( .A(a[3]), .B(b[3]), .Z(n315) );
  GTECH_MUX2 U169 ( .A(n321), .B(n322), .S(n323), .Z(sum[2]) );
  GTECH_NOT U170 ( .A(cin), .Z(n323) );
  GTECH_MUX2 U171 ( .A(n324), .B(n325), .S(n319), .Z(n322) );
  GTECH_OAI21 U172 ( .A(n326), .B(n327), .C(n328), .Z(n319) );
  GTECH_MUX2 U173 ( .A(n325), .B(n324), .S(n329), .Z(n321) );
  GTECH_OAI21 U174 ( .A(b[2]), .B(a[2]), .C(n320), .Z(n324) );
  GTECH_XOR2 U175 ( .A(a[2]), .B(b[2]), .Z(n325) );
  GTECH_MUX2 U176 ( .A(n330), .B(n331), .S(n332), .Z(sum[1]) );
  GTECH_AND_NOT U177 ( .A(n328), .B(n326), .Z(n332) );
  GTECH_OAI21 U178 ( .A(cin), .B(n327), .C(n333), .Z(n331) );
  GTECH_AO21 U179 ( .A(n333), .B(cin), .C(n327), .Z(n330) );
  GTECH_MUX2 U180 ( .A(n334), .B(n335), .S(n336), .Z(sum[15]) );
  GTECH_XOR2 U181 ( .A(n337), .B(n338), .Z(n335) );
  GTECH_OA21 U182 ( .A(n339), .B(n340), .C(n341), .Z(n338) );
  GTECH_XNOR2 U183 ( .A(n337), .B(n342), .Z(n334) );
  GTECH_XNOR2 U184 ( .A(a[15]), .B(b[15]), .Z(n337) );
  GTECH_MUX2 U185 ( .A(n343), .B(n344), .S(n345), .Z(sum[14]) );
  GTECH_OA21 U186 ( .A(n336), .B(n346), .C(n340), .Z(n345) );
  GTECH_OAI21 U187 ( .A(n347), .B(n348), .C(n349), .Z(n340) );
  GTECH_XOR2 U188 ( .A(b[14]), .B(a[14]), .Z(n344) );
  GTECH_OR_NOT U189 ( .A(n339), .B(n341), .Z(n343) );
  GTECH_MUX2 U190 ( .A(n350), .B(n351), .S(n352), .Z(sum[13]) );
  GTECH_MUX2 U191 ( .A(n353), .B(n354), .S(n355), .Z(n351) );
  GTECH_MUX2 U192 ( .A(n353), .B(n354), .S(n347), .Z(n350) );
  GTECH_OR_NOT U193 ( .A(n348), .B(n349), .Z(n354) );
  GTECH_XOR2 U194 ( .A(a[13]), .B(b[13]), .Z(n353) );
  GTECH_XOR2 U195 ( .A(n356), .B(n352), .Z(sum[12]) );
  GTECH_NOT U196 ( .A(n336), .Z(n352) );
  GTECH_MUX2 U197 ( .A(n357), .B(n358), .S(n282), .Z(sum[11]) );
  GTECH_XNOR2 U198 ( .A(n359), .B(n360), .Z(n358) );
  GTECH_AOI21 U199 ( .A(n361), .B(n362), .C(n363), .Z(n360) );
  GTECH_OR2 U200 ( .A(b[10]), .B(a[10]), .Z(n361) );
  GTECH_XOR2 U201 ( .A(n359), .B(n364), .Z(n357) );
  GTECH_XOR2 U202 ( .A(a[11]), .B(b[11]), .Z(n359) );
  GTECH_OAI21 U203 ( .A(n365), .B(n366), .C(n367), .Z(sum[10]) );
  GTECH_MUX2 U204 ( .A(n368), .B(n369), .S(b[10]), .Z(n367) );
  GTECH_OR_NOT U205 ( .A(a[10]), .B(n365), .Z(n369) );
  GTECH_XOR2 U206 ( .A(a[10]), .B(n365), .Z(n368) );
  GTECH_NOT U207 ( .A(n363), .Z(n366) );
  GTECH_AOI21 U208 ( .A(n370), .B(n371), .C(n362), .Z(n365) );
  GTECH_AOI21 U209 ( .A(n281), .B(n285), .C(n284), .Z(n362) );
  GTECH_NOT U210 ( .A(n372), .Z(n284) );
  GTECH_NOT U211 ( .A(n373), .Z(n281) );
  GTECH_XNOR2 U212 ( .A(cin), .B(n374), .Z(sum[0]) );
  GTECH_MUX2 U213 ( .A(n375), .B(n356), .S(n336), .Z(cout) );
  GTECH_OA21 U214 ( .A(n376), .B(n282), .C(n287), .Z(n336) );
  GTECH_OR3 U215 ( .A(n373), .B(n283), .C(n370), .Z(n287) );
  GTECH_NOT U216 ( .A(n288), .Z(n283) );
  GTECH_ADD_AB U217 ( .A(b[8]), .B(a[8]), .COUT(n373) );
  GTECH_NOT U218 ( .A(n370), .Z(n282) );
  GTECH_MUX2 U219 ( .A(n311), .B(n377), .S(n291), .Z(n370) );
  GTECH_NOT U220 ( .A(n312), .Z(n291) );
  GTECH_MUX2 U221 ( .A(n374), .B(n378), .S(cin), .Z(n312) );
  GTECH_AOI21 U222 ( .A(n316), .B(a[3]), .C(n379), .Z(n378) );
  GTECH_OA21 U223 ( .A(a[3]), .B(n316), .C(b[3]), .Z(n379) );
  GTECH_NAND2 U224 ( .A(n380), .B(n320), .Z(n316) );
  GTECH_NAND2 U225 ( .A(a[2]), .B(b[2]), .Z(n320) );
  GTECH_OAI21 U226 ( .A(a[2]), .B(b[2]), .C(n329), .Z(n380) );
  GTECH_OA21 U227 ( .A(n326), .B(n333), .C(n328), .Z(n329) );
  GTECH_OR2 U228 ( .A(b[1]), .B(a[1]), .Z(n328) );
  GTECH_ADD_AB U229 ( .A(b[1]), .B(a[1]), .COUT(n326) );
  GTECH_OR_NOT U230 ( .A(n327), .B(n333), .Z(n374) );
  GTECH_OR2 U231 ( .A(b[0]), .B(a[0]), .Z(n333) );
  GTECH_ADD_AB U232 ( .A(a[0]), .B(b[0]), .COUT(n327) );
  GTECH_OA21 U233 ( .A(a[7]), .B(n293), .C(n381), .Z(n377) );
  GTECH_AO21 U234 ( .A(n293), .B(a[7]), .C(b[7]), .Z(n381) );
  GTECH_NAND2 U235 ( .A(n382), .B(n297), .Z(n293) );
  GTECH_NAND2 U236 ( .A(a[6]), .B(b[6]), .Z(n297) );
  GTECH_OAI21 U237 ( .A(a[6]), .B(b[6]), .C(n302), .Z(n382) );
  GTECH_OA21 U238 ( .A(n305), .B(n310), .C(n306), .Z(n302) );
  GTECH_OR2 U239 ( .A(b[5]), .B(a[5]), .Z(n306) );
  GTECH_ADD_AB U240 ( .A(b[5]), .B(a[5]), .COUT(n305) );
  GTECH_AND_NOT U241 ( .A(n310), .B(n304), .Z(n311) );
  GTECH_ADD_AB U242 ( .A(b[4]), .B(a[4]), .COUT(n304) );
  GTECH_OR2 U243 ( .A(a[4]), .B(b[4]), .Z(n310) );
  GTECH_AOI21 U244 ( .A(n364), .B(a[11]), .C(n383), .Z(n376) );
  GTECH_OA21 U245 ( .A(a[11]), .B(n364), .C(b[11]), .Z(n383) );
  GTECH_OR_NOT U246 ( .A(n363), .B(n384), .Z(n364) );
  GTECH_OAI21 U247 ( .A(a[10]), .B(b[10]), .C(n371), .Z(n384) );
  GTECH_OA21 U248 ( .A(n385), .B(n288), .C(n372), .Z(n371) );
  GTECH_OR2 U249 ( .A(a[9]), .B(b[9]), .Z(n372) );
  GTECH_OR2 U250 ( .A(a[8]), .B(b[8]), .Z(n288) );
  GTECH_NOT U251 ( .A(n285), .Z(n385) );
  GTECH_NAND2 U252 ( .A(b[9]), .B(a[9]), .Z(n285) );
  GTECH_ADD_AB U253 ( .A(a[10]), .B(b[10]), .COUT(n363) );
  GTECH_AND_NOT U254 ( .A(n355), .B(n347), .Z(n356) );
  GTECH_ADD_AB U255 ( .A(b[12]), .B(a[12]), .COUT(n347) );
  GTECH_AO21 U256 ( .A(n342), .B(a[15]), .C(n386), .Z(n375) );
  GTECH_OA21 U257 ( .A(a[15]), .B(n342), .C(b[15]), .Z(n386) );
  GTECH_OAI21 U258 ( .A(n339), .B(n346), .C(n341), .Z(n342) );
  GTECH_OR_NOT U259 ( .A(n387), .B(b[14]), .Z(n341) );
  GTECH_NOT U260 ( .A(a[14]), .Z(n387) );
  GTECH_OAI21 U261 ( .A(n348), .B(n355), .C(n349), .Z(n346) );
  GTECH_OR2 U262 ( .A(a[13]), .B(b[13]), .Z(n349) );
  GTECH_OR2 U263 ( .A(a[12]), .B(b[12]), .Z(n355) );
  GTECH_ADD_AB U264 ( .A(a[13]), .B(b[13]), .COUT(n348) );
  GTECH_NOR2 U265 ( .A(a[14]), .B(b[14]), .Z(n339) );
endmodule

