
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n112, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n112), .K(n112), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n249) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n112), .K(n112), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n112), .K(n112), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n112), .K(n112), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n112), .K(n112), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n112), .K(n112), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]) );
  GTECH_FJK1S A_reg_15_ ( .J(n112), .K(n112), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n265) );
  GTECH_FJK1S A_reg_14_ ( .J(n112), .K(n112), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n264) );
  GTECH_FJK1S A_reg_13_ ( .J(n112), .K(n112), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n263) );
  GTECH_FJK1S A_reg_12_ ( .J(n112), .K(n112), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n262) );
  GTECH_FJK1S A_reg_11_ ( .J(n112), .K(n112), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n261) );
  GTECH_FJK1S A_reg_10_ ( .J(n112), .K(n112), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n260) );
  GTECH_FJK1S A_reg_9_ ( .J(n112), .K(n112), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n259) );
  GTECH_FJK1S A_reg_8_ ( .J(n112), .K(n112), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n258) );
  GTECH_FJK1S A_reg_7_ ( .J(n112), .K(n112), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n257) );
  GTECH_FJK1S A_reg_6_ ( .J(n112), .K(n112), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n256) );
  GTECH_FJK1S A_reg_5_ ( .J(n112), .K(n112), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n255) );
  GTECH_FJK1S A_reg_4_ ( .J(n112), .K(n112), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n254) );
  GTECH_FJK1S A_reg_3_ ( .J(n112), .K(n112), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n253) );
  GTECH_FJK1S A_reg_2_ ( .J(n112), .K(n112), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n252) );
  GTECH_FJK1S A_reg_1_ ( .J(n112), .K(n112), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n251) );
  GTECH_FJK1S A_reg_0_ ( .J(n112), .K(n112), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n250) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n112), .K(n112), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n112), .K(n112), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n112), .K(n112), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n112), .K(n112), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n112), .K(n112), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n112), .K(n112), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n112), .K(n112), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n112), .K(n112), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n112), .K(n112), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n112), .K(n112), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n112), .K(n112), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n112), .K(n112), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n112), .K(n112), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n112), .K(n112), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n112), .K(n112), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n112), .K(n112), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n112), .K(n112), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n112), .K(n112), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n112), .K(n112), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n112), .K(n112), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n112), .K(n112), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n112), .K(n112), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n112), .K(n112), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n112), .K(n112), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n112), .K(n112), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n112), .K(n112), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n112), .K(n112), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n112), .K(n112), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n112), .K(n112), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n112), .K(n112), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n112), .K(n112), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n112), .K(n112), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n112), .K(n112), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n112), .K(n112), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n112), .K(n112), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n112), .K(n112), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n112), .K(n112), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n112), .K(n112), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n112), .K(n112), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n112), .K(n112), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n112), .K(n112), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n112), .K(n112), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n112), .K(n112), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n112), .K(n112), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n112), .K(n112), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n112), .K(n112), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n112), .K(n112), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n112), .K(n112), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n112), .K(n112), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n112), .K(n112), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n112), .K(n112), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n112), .K(n112), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n112), .K(n112), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n112), .K(n112), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n112), .K(n112), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n112), .K(n112), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n112), .K(n112), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n112), .K(n112), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n112), .K(n112), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n112), .K(n112), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n112), .K(n112), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n112), .K(n112), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n112), .K(n112), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n112), .K(n112), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n112), .K(n112), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n112), .K(n112), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U251 ( .Z(n112) );
  GTECH_NOT U252 ( .A(n267), .Z(N99) );
  GTECH_AOI222 U253 ( .A(n268), .B(n269), .C(n270), .D(n271), .E(n272), .F(
        n273), .Z(n267) );
  GTECH_NOT U254 ( .A(n274), .Z(N98) );
  GTECH_AOI222 U255 ( .A(n270), .B(n275), .C(n276), .D(n277), .E(R[15]), .F(
        n278), .Z(n274) );
  GTECH_NAND2 U256 ( .A(n279), .B(n280), .Z(n276) );
  GTECH_OAI2N2 U257 ( .A(n13), .B(n281), .C(R[14]), .D(n278), .Z(N97) );
  GTECH_OAI2N2 U258 ( .A(n14), .B(n281), .C(R[13]), .D(n278), .Z(N96) );
  GTECH_OAI2N2 U259 ( .A(n15), .B(n281), .C(R[12]), .D(n278), .Z(N95) );
  GTECH_OAI2N2 U260 ( .A(n16), .B(n281), .C(R[11]), .D(n278), .Z(N94) );
  GTECH_OAI2N2 U261 ( .A(n17), .B(n281), .C(R[10]), .D(n278), .Z(N93) );
  GTECH_OAI2N2 U262 ( .A(n18), .B(n281), .C(R[9]), .D(n278), .Z(N92) );
  GTECH_OAI2N2 U263 ( .A(n19), .B(n281), .C(R[8]), .D(n278), .Z(N91) );
  GTECH_OAI2N2 U264 ( .A(n20), .B(n281), .C(R[7]), .D(n278), .Z(N90) );
  GTECH_OAI2N2 U265 ( .A(n21), .B(n281), .C(R[6]), .D(n278), .Z(N89) );
  GTECH_OAI2N2 U266 ( .A(n22), .B(n281), .C(R[5]), .D(n278), .Z(N88) );
  GTECH_OAI2N2 U267 ( .A(n23), .B(n281), .C(R[4]), .D(n278), .Z(N87) );
  GTECH_OAI2N2 U268 ( .A(n24), .B(n281), .C(R[3]), .D(n278), .Z(N86) );
  GTECH_OAI2N2 U269 ( .A(n25), .B(n281), .C(R[2]), .D(n278), .Z(N85) );
  GTECH_OAI2N2 U270 ( .A(n26), .B(n281), .C(R[1]), .D(n278), .Z(N84) );
  GTECH_OAI2N2 U271 ( .A(n27), .B(n281), .C(R[0]), .D(n278), .Z(N83) );
  GTECH_AND2 U272 ( .A(M[15]), .B(n278), .Z(N42) );
  GTECH_AND2 U273 ( .A(M[14]), .B(n278), .Z(N39) );
  GTECH_AND2 U274 ( .A(M[13]), .B(n278), .Z(N38) );
  GTECH_AND2 U275 ( .A(M[12]), .B(n278), .Z(N37) );
  GTECH_AND2 U276 ( .A(M[11]), .B(n278), .Z(N36) );
  GTECH_AND2 U277 ( .A(M[10]), .B(n278), .Z(N35) );
  GTECH_AND2 U278 ( .A(M[9]), .B(n278), .Z(N34) );
  GTECH_AND2 U279 ( .A(M[8]), .B(n278), .Z(N33) );
  GTECH_AND2 U280 ( .A(M[7]), .B(n278), .Z(N32) );
  GTECH_AND2 U281 ( .A(M[6]), .B(n278), .Z(N31) );
  GTECH_AND2 U282 ( .A(M[5]), .B(n278), .Z(N30) );
  GTECH_AND2 U283 ( .A(M[4]), .B(n278), .Z(N29) );
  GTECH_AND2 U284 ( .A(M[3]), .B(n278), .Z(N28) );
  GTECH_AND2 U285 ( .A(M[2]), .B(n278), .Z(N27) );
  GTECH_AND2 U286 ( .A(M[1]), .B(n278), .Z(N26) );
  GTECH_AND2 U287 ( .A(M[0]), .B(n278), .Z(N25) );
  GTECH_NOT U288 ( .A(n282), .Z(n278) );
  GTECH_OAI21 U289 ( .A(n9), .B(n283), .C(n282), .Z(N19) );
  GTECH_OR_NOT U290 ( .A(n281), .B(n284), .Z(n283) );
  GTECH_OR3 U291 ( .A(Rst), .B(Ld), .C(n285), .Z(N18) );
  GTECH_AND2 U292 ( .A(n285), .B(n286), .Z(N17) );
  GTECH_OAI21 U293 ( .A(n8), .B(n287), .C(n284), .Z(n286) );
  GTECH_AND2 U294 ( .A(n285), .B(n288), .Z(N16) );
  GTECH_OAI21 U295 ( .A(n7), .B(n289), .C(n290), .Z(n288) );
  GTECH_NOT U296 ( .A(n291), .Z(N152) );
  GTECH_AOI222 U297 ( .A(n292), .B(n293), .C(n294), .D(n295), .E(n296), .F(
        n297), .Z(n291) );
  GTECH_NAND2 U298 ( .A(n298), .B(n299), .Z(N151) );
  GTECH_NOT U299 ( .A(n300), .Z(N150) );
  GTECH_AOI222 U300 ( .A(n301), .B(n292), .C(n294), .D(n302), .E(n296), .F(
        n303), .Z(n300) );
  GTECH_MUX2 U301 ( .A(n304), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND_NOT U302 ( .A(n285), .B(n249), .Z(n304) );
  GTECH_NOT U303 ( .A(n305), .Z(N149) );
  GTECH_AOI222 U304 ( .A(n306), .B(n292), .C(n294), .D(n307), .E(n296), .F(
        n308), .Z(n305) );
  GTECH_NOT U305 ( .A(n309), .Z(N148) );
  GTECH_AOI222 U306 ( .A(n310), .B(n292), .C(n294), .D(n311), .E(n296), .F(
        n312), .Z(n309) );
  GTECH_NOT U307 ( .A(n313), .Z(N147) );
  GTECH_AOI222 U308 ( .A(n314), .B(n292), .C(n294), .D(n315), .E(n296), .F(
        n316), .Z(n313) );
  GTECH_NOT U309 ( .A(n317), .Z(N146) );
  GTECH_AOI222 U310 ( .A(n318), .B(n292), .C(n294), .D(n319), .E(n296), .F(
        n320), .Z(n317) );
  GTECH_NOT U311 ( .A(n321), .Z(N145) );
  GTECH_AOI222 U312 ( .A(n322), .B(n292), .C(n294), .D(n323), .E(n296), .F(
        n324), .Z(n321) );
  GTECH_NOT U313 ( .A(n325), .Z(N144) );
  GTECH_AOI222 U314 ( .A(n326), .B(n292), .C(n294), .D(n327), .E(n296), .F(
        n328), .Z(n325) );
  GTECH_NOT U315 ( .A(n329), .Z(N143) );
  GTECH_AOI222 U316 ( .A(n330), .B(n292), .C(n294), .D(n331), .E(n296), .F(
        n332), .Z(n329) );
  GTECH_NOT U317 ( .A(n333), .Z(N142) );
  GTECH_AOI222 U318 ( .A(n334), .B(n292), .C(n294), .D(n335), .E(n296), .F(
        n336), .Z(n333) );
  GTECH_NOT U319 ( .A(n337), .Z(N141) );
  GTECH_AOI222 U320 ( .A(n338), .B(n292), .C(n294), .D(n339), .E(n296), .F(
        n340), .Z(n337) );
  GTECH_NOT U321 ( .A(n341), .Z(N140) );
  GTECH_AOI222 U322 ( .A(n342), .B(n292), .C(n294), .D(n343), .E(n296), .F(
        n344), .Z(n341) );
  GTECH_NOT U323 ( .A(n345), .Z(N14) );
  GTECH_NAND2 U324 ( .A(n285), .B(n249), .Z(n345) );
  GTECH_NOT U325 ( .A(n346), .Z(N139) );
  GTECH_AOI222 U326 ( .A(n347), .B(n292), .C(n294), .D(n348), .E(n296), .F(
        n349), .Z(n346) );
  GTECH_NOT U327 ( .A(n350), .Z(N138) );
  GTECH_AOI222 U328 ( .A(n351), .B(n292), .C(n294), .D(n352), .E(n296), .F(
        n353), .Z(n350) );
  GTECH_NOT U329 ( .A(n354), .Z(N137) );
  GTECH_AOI222 U330 ( .A(n355), .B(n292), .C(n294), .D(n356), .E(n296), .F(
        n357), .Z(n354) );
  GTECH_NOT U331 ( .A(n358), .Z(N136) );
  GTECH_AOI222 U332 ( .A(n292), .B(n269), .C(n294), .D(n271), .E(n296), .F(
        n273), .Z(n358) );
  GTECH_NOT U333 ( .A(n359), .Z(n273) );
  GTECH_XOR2 U334 ( .A(n360), .B(n361), .Z(n359) );
  GTECH_NOT U335 ( .A(n362), .Z(n361) );
  GTECH_NOT U336 ( .A(n363), .Z(n294) );
  GTECH_NOT U337 ( .A(n364), .Z(n269) );
  GTECH_XOR2 U338 ( .A(n360), .B(n365), .Z(n364) );
  GTECH_NOT U339 ( .A(n366), .Z(n365) );
  GTECH_XOR2 U340 ( .A(n271), .B(n251), .Z(n360) );
  GTECH_OAI21 U341 ( .A(n12), .B(n363), .C(n367), .Z(N135) );
  GTECH_OAI21 U342 ( .A(n296), .B(n292), .C(n277), .Z(n367) );
  GTECH_OAI21 U343 ( .A(n12), .B(n368), .C(n362), .Z(n277) );
  GTECH_NOT U344 ( .A(n369), .Z(n292) );
  GTECH_OR3 U345 ( .A(n10), .B(n370), .C(n299), .Z(n369) );
  GTECH_NOT U346 ( .A(n371), .Z(n296) );
  GTECH_OR3 U347 ( .A(n28), .B(n372), .C(n299), .Z(n371) );
  GTECH_NAND2 U348 ( .A(n373), .B(N155), .Z(n363) );
  GTECH_XOR2 U349 ( .A(n372), .B(n28), .Z(n373) );
  GTECH_NOT U350 ( .A(n10), .Z(n372) );
  GTECH_AND2 U351 ( .A(N155), .B(n374), .Z(N134) );
  GTECH_NOT U352 ( .A(n13), .Z(n374) );
  GTECH_AND2 U353 ( .A(N155), .B(n375), .Z(N133) );
  GTECH_NOT U354 ( .A(n14), .Z(n375) );
  GTECH_AND2 U355 ( .A(N155), .B(n376), .Z(N132) );
  GTECH_NOT U356 ( .A(n15), .Z(n376) );
  GTECH_AND2 U357 ( .A(N155), .B(n377), .Z(N131) );
  GTECH_NOT U358 ( .A(n16), .Z(n377) );
  GTECH_AND2 U359 ( .A(N155), .B(n378), .Z(N130) );
  GTECH_NOT U360 ( .A(n17), .Z(n378) );
  GTECH_AND2 U361 ( .A(N155), .B(n379), .Z(N129) );
  GTECH_NOT U362 ( .A(n18), .Z(n379) );
  GTECH_AND2 U363 ( .A(N155), .B(n380), .Z(N128) );
  GTECH_NOT U364 ( .A(n19), .Z(n380) );
  GTECH_AND2 U365 ( .A(N155), .B(n381), .Z(N127) );
  GTECH_NOT U366 ( .A(n20), .Z(n381) );
  GTECH_AND2 U367 ( .A(N155), .B(n382), .Z(N126) );
  GTECH_NOT U368 ( .A(n21), .Z(n382) );
  GTECH_AND2 U369 ( .A(N155), .B(n383), .Z(N125) );
  GTECH_NOT U370 ( .A(n22), .Z(n383) );
  GTECH_AND2 U371 ( .A(N155), .B(n384), .Z(N124) );
  GTECH_NOT U372 ( .A(n23), .Z(n384) );
  GTECH_AND2 U373 ( .A(N155), .B(n385), .Z(N123) );
  GTECH_NOT U374 ( .A(n24), .Z(n385) );
  GTECH_AND2 U375 ( .A(N155), .B(n386), .Z(N122) );
  GTECH_NOT U376 ( .A(n25), .Z(n386) );
  GTECH_AND2 U377 ( .A(N155), .B(n387), .Z(N121) );
  GTECH_NOT U378 ( .A(n26), .Z(n387) );
  GTECH_AND2 U379 ( .A(N155), .B(n388), .Z(N120) );
  GTECH_NOT U380 ( .A(n27), .Z(n388) );
  GTECH_NOT U381 ( .A(n299), .Z(N155) );
  GTECH_NAND5 U382 ( .A(n389), .B(n6), .C(n9), .D(n8), .E(n7), .Z(n299) );
  GTECH_NOR2 U383 ( .A(n249), .B(Rst), .Z(n389) );
  GTECH_NOT U384 ( .A(n390), .Z(N116) );
  GTECH_AOI222 U385 ( .A(n270), .B(n295), .C(n272), .D(n297), .E(n293), .F(
        n268), .Z(n390) );
  GTECH_XOR2 U386 ( .A(n391), .B(n392), .Z(n293) );
  GTECH_ADD_ABC U387 ( .A(n31), .B(n265), .C(n393), .COUT(n392) );
  GTECH_XOR2 U388 ( .A(n394), .B(n391), .Z(n297) );
  GTECH_XOR2 U389 ( .A(A[16]), .B(n30), .Z(n391) );
  GTECH_OAI21 U390 ( .A(n395), .B(n31), .C(n396), .Z(n394) );
  GTECH_OAI21 U391 ( .A(n265), .B(n302), .C(n397), .Z(n396) );
  GTECH_NOT U392 ( .A(n30), .Z(n295) );
  GTECH_NAND2 U393 ( .A(n281), .B(n398), .Z(N115) );
  GTECH_NOT U394 ( .A(N41), .Z(n398) );
  GTECH_NAND2 U395 ( .A(n298), .B(n282), .Z(N41) );
  GTECH_NAND2 U396 ( .A(Ld), .B(n298), .Z(n282) );
  GTECH_NOT U397 ( .A(Rst), .Z(n298) );
  GTECH_NOT U398 ( .A(n399), .Z(N113) );
  GTECH_AOI222 U399 ( .A(n270), .B(n302), .C(n272), .D(n303), .E(n301), .F(
        n268), .Z(n399) );
  GTECH_XOR2 U400 ( .A(n400), .B(n393), .Z(n301) );
  GTECH_ADD_ABC U401 ( .A(n32), .B(n264), .C(n401), .COUT(n393) );
  GTECH_NOT U402 ( .A(n402), .Z(n303) );
  GTECH_XOR2 U403 ( .A(n400), .B(n403), .Z(n402) );
  GTECH_NOT U404 ( .A(n397), .Z(n403) );
  GTECH_OAI21 U405 ( .A(n32), .B(n404), .C(n405), .Z(n397) );
  GTECH_OAI21 U406 ( .A(n264), .B(n307), .C(n406), .Z(n405) );
  GTECH_XOR2 U407 ( .A(n395), .B(n31), .Z(n400) );
  GTECH_NOT U408 ( .A(n265), .Z(n395) );
  GTECH_NOT U409 ( .A(n31), .Z(n302) );
  GTECH_NOT U410 ( .A(n407), .Z(N112) );
  GTECH_AOI222 U411 ( .A(n270), .B(n307), .C(n272), .D(n308), .E(n306), .F(
        n268), .Z(n407) );
  GTECH_XOR2 U412 ( .A(n408), .B(n401), .Z(n306) );
  GTECH_ADD_ABC U413 ( .A(n33), .B(n263), .C(n409), .COUT(n401) );
  GTECH_NOT U414 ( .A(n410), .Z(n308) );
  GTECH_XOR2 U415 ( .A(n408), .B(n411), .Z(n410) );
  GTECH_NOT U416 ( .A(n406), .Z(n411) );
  GTECH_OAI21 U417 ( .A(n33), .B(n412), .C(n413), .Z(n406) );
  GTECH_OAI21 U418 ( .A(n263), .B(n311), .C(n414), .Z(n413) );
  GTECH_XOR2 U419 ( .A(n404), .B(n32), .Z(n408) );
  GTECH_NOT U420 ( .A(n264), .Z(n404) );
  GTECH_NOT U421 ( .A(n32), .Z(n307) );
  GTECH_NOT U422 ( .A(n415), .Z(N111) );
  GTECH_AOI222 U423 ( .A(n270), .B(n311), .C(n272), .D(n312), .E(n310), .F(
        n268), .Z(n415) );
  GTECH_XOR2 U424 ( .A(n416), .B(n409), .Z(n310) );
  GTECH_ADD_ABC U425 ( .A(n34), .B(n262), .C(n417), .COUT(n409) );
  GTECH_NOT U426 ( .A(n418), .Z(n312) );
  GTECH_XOR2 U427 ( .A(n416), .B(n419), .Z(n418) );
  GTECH_NOT U428 ( .A(n414), .Z(n419) );
  GTECH_OAI21 U429 ( .A(n34), .B(n420), .C(n421), .Z(n414) );
  GTECH_OAI21 U430 ( .A(n262), .B(n315), .C(n422), .Z(n421) );
  GTECH_XOR2 U431 ( .A(n412), .B(n33), .Z(n416) );
  GTECH_NOT U432 ( .A(n263), .Z(n412) );
  GTECH_NOT U433 ( .A(n33), .Z(n311) );
  GTECH_NOT U434 ( .A(n423), .Z(N110) );
  GTECH_AOI222 U435 ( .A(n270), .B(n315), .C(n272), .D(n316), .E(n314), .F(
        n268), .Z(n423) );
  GTECH_XOR2 U436 ( .A(n424), .B(n417), .Z(n314) );
  GTECH_ADD_ABC U437 ( .A(n35), .B(n261), .C(n425), .COUT(n417) );
  GTECH_NOT U438 ( .A(n426), .Z(n316) );
  GTECH_XOR2 U439 ( .A(n424), .B(n427), .Z(n426) );
  GTECH_NOT U440 ( .A(n422), .Z(n427) );
  GTECH_OAI21 U441 ( .A(n35), .B(n428), .C(n429), .Z(n422) );
  GTECH_OAI21 U442 ( .A(n261), .B(n319), .C(n430), .Z(n429) );
  GTECH_XOR2 U443 ( .A(n420), .B(n34), .Z(n424) );
  GTECH_NOT U444 ( .A(n262), .Z(n420) );
  GTECH_NOT U445 ( .A(n34), .Z(n315) );
  GTECH_NOT U446 ( .A(n431), .Z(N109) );
  GTECH_AOI222 U447 ( .A(n270), .B(n319), .C(n272), .D(n320), .E(n318), .F(
        n268), .Z(n431) );
  GTECH_XOR2 U448 ( .A(n432), .B(n425), .Z(n318) );
  GTECH_ADD_ABC U449 ( .A(n36), .B(n260), .C(n433), .COUT(n425) );
  GTECH_NOT U450 ( .A(n434), .Z(n320) );
  GTECH_XOR2 U451 ( .A(n432), .B(n435), .Z(n434) );
  GTECH_NOT U452 ( .A(n430), .Z(n435) );
  GTECH_OAI21 U453 ( .A(n36), .B(n436), .C(n437), .Z(n430) );
  GTECH_OAI21 U454 ( .A(n260), .B(n323), .C(n438), .Z(n437) );
  GTECH_XOR2 U455 ( .A(n428), .B(n35), .Z(n432) );
  GTECH_NOT U456 ( .A(n261), .Z(n428) );
  GTECH_NOT U457 ( .A(n35), .Z(n319) );
  GTECH_NOT U458 ( .A(n439), .Z(N108) );
  GTECH_AOI222 U459 ( .A(n270), .B(n323), .C(n272), .D(n324), .E(n322), .F(
        n268), .Z(n439) );
  GTECH_XOR2 U460 ( .A(n440), .B(n433), .Z(n322) );
  GTECH_ADD_ABC U461 ( .A(n37), .B(n259), .C(n441), .COUT(n433) );
  GTECH_NOT U462 ( .A(n442), .Z(n324) );
  GTECH_XOR2 U463 ( .A(n440), .B(n443), .Z(n442) );
  GTECH_NOT U464 ( .A(n438), .Z(n443) );
  GTECH_OAI21 U465 ( .A(n37), .B(n444), .C(n445), .Z(n438) );
  GTECH_OAI21 U466 ( .A(n259), .B(n327), .C(n446), .Z(n445) );
  GTECH_XOR2 U467 ( .A(n436), .B(n36), .Z(n440) );
  GTECH_NOT U468 ( .A(n260), .Z(n436) );
  GTECH_NOT U469 ( .A(n36), .Z(n323) );
  GTECH_NOT U470 ( .A(n447), .Z(N107) );
  GTECH_AOI222 U471 ( .A(n270), .B(n327), .C(n272), .D(n328), .E(n326), .F(
        n268), .Z(n447) );
  GTECH_XOR2 U472 ( .A(n448), .B(n441), .Z(n326) );
  GTECH_ADD_ABC U473 ( .A(n38), .B(n258), .C(n449), .COUT(n441) );
  GTECH_NOT U474 ( .A(n450), .Z(n328) );
  GTECH_XOR2 U475 ( .A(n448), .B(n451), .Z(n450) );
  GTECH_NOT U476 ( .A(n446), .Z(n451) );
  GTECH_OAI21 U477 ( .A(n38), .B(n452), .C(n453), .Z(n446) );
  GTECH_OAI21 U478 ( .A(n258), .B(n331), .C(n454), .Z(n453) );
  GTECH_XOR2 U479 ( .A(n444), .B(n37), .Z(n448) );
  GTECH_NOT U480 ( .A(n259), .Z(n444) );
  GTECH_NOT U481 ( .A(n37), .Z(n327) );
  GTECH_NOT U482 ( .A(n455), .Z(N106) );
  GTECH_AOI222 U483 ( .A(n270), .B(n331), .C(n272), .D(n332), .E(n330), .F(
        n268), .Z(n455) );
  GTECH_XOR2 U484 ( .A(n456), .B(n449), .Z(n330) );
  GTECH_ADD_ABC U485 ( .A(n39), .B(n257), .C(n457), .COUT(n449) );
  GTECH_NOT U486 ( .A(n458), .Z(n332) );
  GTECH_XOR2 U487 ( .A(n456), .B(n459), .Z(n458) );
  GTECH_NOT U488 ( .A(n454), .Z(n459) );
  GTECH_OAI21 U489 ( .A(n39), .B(n460), .C(n461), .Z(n454) );
  GTECH_OAI21 U490 ( .A(n257), .B(n335), .C(n462), .Z(n461) );
  GTECH_XOR2 U491 ( .A(n452), .B(n38), .Z(n456) );
  GTECH_NOT U492 ( .A(n258), .Z(n452) );
  GTECH_NOT U493 ( .A(n38), .Z(n331) );
  GTECH_NOT U494 ( .A(n463), .Z(N105) );
  GTECH_AOI222 U495 ( .A(n270), .B(n335), .C(n272), .D(n336), .E(n334), .F(
        n268), .Z(n463) );
  GTECH_XOR2 U496 ( .A(n464), .B(n457), .Z(n334) );
  GTECH_ADD_ABC U497 ( .A(n40), .B(n256), .C(n465), .COUT(n457) );
  GTECH_NOT U498 ( .A(n466), .Z(n336) );
  GTECH_XOR2 U499 ( .A(n464), .B(n467), .Z(n466) );
  GTECH_NOT U500 ( .A(n462), .Z(n467) );
  GTECH_OAI21 U501 ( .A(n40), .B(n468), .C(n469), .Z(n462) );
  GTECH_OAI21 U502 ( .A(n256), .B(n339), .C(n470), .Z(n469) );
  GTECH_XOR2 U503 ( .A(n460), .B(n39), .Z(n464) );
  GTECH_NOT U504 ( .A(n257), .Z(n460) );
  GTECH_NOT U505 ( .A(n39), .Z(n335) );
  GTECH_NOT U506 ( .A(n471), .Z(N104) );
  GTECH_AOI222 U507 ( .A(n270), .B(n339), .C(n272), .D(n340), .E(n338), .F(
        n268), .Z(n471) );
  GTECH_XOR2 U508 ( .A(n472), .B(n465), .Z(n338) );
  GTECH_ADD_ABC U509 ( .A(n41), .B(n255), .C(n473), .COUT(n465) );
  GTECH_NOT U510 ( .A(n474), .Z(n340) );
  GTECH_XOR2 U511 ( .A(n472), .B(n475), .Z(n474) );
  GTECH_NOT U512 ( .A(n470), .Z(n475) );
  GTECH_OAI21 U513 ( .A(n41), .B(n476), .C(n477), .Z(n470) );
  GTECH_OAI21 U514 ( .A(n255), .B(n343), .C(n478), .Z(n477) );
  GTECH_XOR2 U515 ( .A(n468), .B(n40), .Z(n472) );
  GTECH_NOT U516 ( .A(n256), .Z(n468) );
  GTECH_NOT U517 ( .A(n40), .Z(n339) );
  GTECH_NOT U518 ( .A(n479), .Z(N103) );
  GTECH_AOI222 U519 ( .A(n270), .B(n343), .C(n272), .D(n344), .E(n342), .F(
        n268), .Z(n479) );
  GTECH_XOR2 U520 ( .A(n480), .B(n473), .Z(n342) );
  GTECH_ADD_ABC U521 ( .A(n42), .B(n254), .C(n481), .COUT(n473) );
  GTECH_NOT U522 ( .A(n482), .Z(n344) );
  GTECH_XOR2 U523 ( .A(n480), .B(n483), .Z(n482) );
  GTECH_NOT U524 ( .A(n478), .Z(n483) );
  GTECH_OAI21 U525 ( .A(n42), .B(n484), .C(n485), .Z(n478) );
  GTECH_OAI21 U526 ( .A(n254), .B(n348), .C(n486), .Z(n485) );
  GTECH_XOR2 U527 ( .A(n476), .B(n41), .Z(n480) );
  GTECH_NOT U528 ( .A(n255), .Z(n476) );
  GTECH_NOT U529 ( .A(n41), .Z(n343) );
  GTECH_NOT U530 ( .A(n487), .Z(N102) );
  GTECH_AOI222 U531 ( .A(n270), .B(n348), .C(n272), .D(n349), .E(n347), .F(
        n268), .Z(n487) );
  GTECH_XOR2 U532 ( .A(n488), .B(n481), .Z(n347) );
  GTECH_ADD_ABC U533 ( .A(n43), .B(n253), .C(n489), .COUT(n481) );
  GTECH_NOT U534 ( .A(n490), .Z(n349) );
  GTECH_XOR2 U535 ( .A(n488), .B(n491), .Z(n490) );
  GTECH_NOT U536 ( .A(n486), .Z(n491) );
  GTECH_OAI21 U537 ( .A(n43), .B(n492), .C(n493), .Z(n486) );
  GTECH_OAI21 U538 ( .A(n253), .B(n352), .C(n494), .Z(n493) );
  GTECH_XOR2 U539 ( .A(n484), .B(n42), .Z(n488) );
  GTECH_NOT U540 ( .A(n254), .Z(n484) );
  GTECH_NOT U541 ( .A(n42), .Z(n348) );
  GTECH_NOT U542 ( .A(n495), .Z(N101) );
  GTECH_AOI222 U543 ( .A(n270), .B(n352), .C(n272), .D(n353), .E(n351), .F(
        n268), .Z(n495) );
  GTECH_XOR2 U544 ( .A(n496), .B(n489), .Z(n351) );
  GTECH_ADD_ABC U545 ( .A(n29), .B(n252), .C(n497), .COUT(n489) );
  GTECH_NOT U546 ( .A(n498), .Z(n353) );
  GTECH_XOR2 U547 ( .A(n496), .B(n499), .Z(n498) );
  GTECH_NOT U548 ( .A(n494), .Z(n499) );
  GTECH_OAI21 U549 ( .A(n29), .B(n500), .C(n501), .Z(n494) );
  GTECH_OAI21 U550 ( .A(n252), .B(n356), .C(n502), .Z(n501) );
  GTECH_XOR2 U551 ( .A(n492), .B(n43), .Z(n496) );
  GTECH_NOT U552 ( .A(n253), .Z(n492) );
  GTECH_NOT U553 ( .A(n43), .Z(n352) );
  GTECH_NOT U554 ( .A(n503), .Z(N100) );
  GTECH_AOI222 U555 ( .A(n355), .B(n268), .C(n270), .D(n356), .E(n272), .F(
        n357), .Z(n503) );
  GTECH_NOT U556 ( .A(n504), .Z(n357) );
  GTECH_XOR2 U557 ( .A(n505), .B(n506), .Z(n504) );
  GTECH_NOT U558 ( .A(n502), .Z(n506) );
  GTECH_OAI21 U559 ( .A(n11), .B(n507), .C(n508), .Z(n502) );
  GTECH_OAI21 U560 ( .A(n251), .B(n271), .C(n362), .Z(n508) );
  GTECH_NAND2 U561 ( .A(n12), .B(n368), .Z(n362) );
  GTECH_NOT U562 ( .A(n11), .Z(n271) );
  GTECH_NOT U563 ( .A(n251), .Z(n507) );
  GTECH_NOT U564 ( .A(n280), .Z(n272) );
  GTECH_NAND2 U565 ( .A(N82), .B(n10), .Z(n280) );
  GTECH_NOT U566 ( .A(n509), .Z(N82) );
  GTECH_NOT U567 ( .A(n29), .Z(n356) );
  GTECH_NOT U568 ( .A(n510), .Z(n270) );
  GTECH_MUX2 U569 ( .A(n509), .B(n511), .S(n10), .Z(n510) );
  GTECH_NAND2 U570 ( .A(n28), .B(n285), .Z(n511) );
  GTECH_NAND2 U571 ( .A(n285), .B(n370), .Z(n509) );
  GTECH_NOT U572 ( .A(n281), .Z(n285) );
  GTECH_NOT U573 ( .A(n279), .Z(n268) );
  GTECH_OR3 U574 ( .A(n10), .B(n281), .C(n370), .Z(n279) );
  GTECH_NOT U575 ( .A(n28), .Z(n370) );
  GTECH_OR3 U576 ( .A(Ld), .B(Rst), .C(n512), .Z(n281) );
  GTECH_AND_NOT U577 ( .A(n9), .B(n284), .Z(n512) );
  GTECH_NAND2 U578 ( .A(n8), .B(n287), .Z(n284) );
  GTECH_NOT U579 ( .A(n290), .Z(n287) );
  GTECH_NAND2 U580 ( .A(n7), .B(n289), .Z(n290) );
  GTECH_NOT U581 ( .A(n513), .Z(n289) );
  GTECH_NAND2 U582 ( .A(n6), .B(n249), .Z(n513) );
  GTECH_XOR2 U583 ( .A(n505), .B(n497), .Z(n355) );
  GTECH_ADD_ABC U584 ( .A(n251), .B(n11), .C(n366), .COUT(n497) );
  GTECH_NAND2 U585 ( .A(n275), .B(n368), .Z(n366) );
  GTECH_NOT U586 ( .A(n250), .Z(n368) );
  GTECH_NOT U587 ( .A(n12), .Z(n275) );
  GTECH_XOR2 U588 ( .A(n500), .B(n29), .Z(n505) );
  GTECH_NOT U589 ( .A(n252), .Z(n500) );
endmodule

