
module fraction_multiplier4 ( CLK, St, Mplier, Mcand, Product, Done );
  input [3:0] Mplier;
  input [3:0] Mcand;
  output [6:0] Product;
  input CLK, St;
  output Done;
  wire   N40, N41, N42, N44, N46, N48, N50, N52, N54, N56, N57, N58, N63, n12,
         n13, n14, n16, n17, n18, n19, n20, n75, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;
  wire   [2:0] State;

  GTECH_FD1 State_reg_0_ ( .D(N40), .CP(CLK), .Q(State[0]), .QN(n12) );
  GTECH_FD1 State_reg_2_ ( .D(N42), .CP(CLK), .Q(State[2]), .QN(n13) );
  GTECH_FD1 State_reg_1_ ( .D(N41), .CP(CLK), .Q(State[1]), .QN(n85) );
  GTECH_FJK1S B_reg_0_ ( .J(n75), .K(n75), .TI(N52), .TE(N57), .CP(CLK), .Q(
        Product[0]), .QN(n14) );
  GTECH_FJK1S A_reg_3_ ( .J(n75), .K(n75), .TI(N50), .TE(N63), .CP(CLK), .QN(
        n83) );
  GTECH_FJK1S A_reg_0_ ( .J(n75), .K(n75), .TI(N44), .TE(N57), .CP(CLK), .Q(
        Product[4]), .QN(n16) );
  GTECH_FJK1S A_reg_1_ ( .J(n75), .K(n75), .TI(N46), .TE(N57), .CP(CLK), .Q(
        Product[5]), .QN(n17) );
  GTECH_FJK1S A_reg_2_ ( .J(n75), .K(n75), .TI(N48), .TE(N57), .CP(CLK), .Q(
        Product[6]), .QN(n84) );
  GTECH_FJK1S B_reg_3_ ( .J(n75), .K(n75), .TI(N58), .TE(N57), .CP(CLK), .Q(
        Product[3]), .QN(n18) );
  GTECH_FJK1S B_reg_2_ ( .J(n75), .K(n75), .TI(N56), .TE(N57), .CP(CLK), .Q(
        Product[2]), .QN(n19) );
  GTECH_FJK1S B_reg_1_ ( .J(n75), .K(n75), .TI(N54), .TE(N57), .CP(CLK), .Q(
        Product[1]), .QN(n20) );
  GTECH_ZERO U79 ( .Z(n75) );
  GTECH_AND2 U80 ( .A(n86), .B(N57), .Z(N63) );
  GTECH_NOT U81 ( .A(n87), .Z(N58) );
  GTECH_AOI222 U82 ( .A(Mplier[3]), .B(n88), .C(n89), .D(n90), .E(n91), .F(n92), .Z(n87) );
  GTECH_OAI21 U83 ( .A(Mcand[0]), .B(n93), .C(n86), .Z(n91) );
  GTECH_NOR2 U84 ( .A(n14), .B(n93), .Z(n89) );
  GTECH_OAI21 U85 ( .A(n94), .B(n95), .C(n93), .Z(N57) );
  GTECH_OAI2N2 U86 ( .A(n18), .B(n93), .C(Mplier[2]), .D(n88), .Z(N56) );
  GTECH_OAI2N2 U87 ( .A(n19), .B(n93), .C(Mplier[1]), .D(n88), .Z(N54) );
  GTECH_OAI2N2 U88 ( .A(n20), .B(n93), .C(Mplier[0]), .D(n88), .Z(N52) );
  GTECH_MUX2 U89 ( .A(n96), .B(n97), .S(Mcand[3]), .Z(N50) );
  GTECH_MUX2 U90 ( .A(n98), .B(n99), .S(n83), .Z(N48) );
  GTECH_NOT U91 ( .A(n100), .Z(n99) );
  GTECH_MUX2 U92 ( .A(n101), .B(n102), .S(Mcand[3]), .Z(n100) );
  GTECH_NAND2 U93 ( .A(n103), .B(n86), .Z(n98) );
  GTECH_MUX2 U94 ( .A(n102), .B(n101), .S(Mcand[3]), .Z(n103) );
  GTECH_OA22 U95 ( .A(n104), .B(n105), .C(n106), .D(n107), .Z(n101) );
  GTECH_AOI22 U96 ( .A(n104), .B(n108), .C(n106), .D(n109), .Z(n102) );
  GTECH_OA21 U97 ( .A(n110), .B(n111), .C(n112), .Z(n106) );
  GTECH_AO21 U98 ( .A(n110), .B(n111), .C(n84), .Z(n112) );
  GTECH_OA21 U99 ( .A(n111), .B(n113), .C(n114), .Z(n104) );
  GTECH_OAI21 U100 ( .A(n115), .B(Mcand[2]), .C(n84), .Z(n114) );
  GTECH_MUX2 U101 ( .A(n116), .B(n117), .S(n84), .Z(N46) );
  GTECH_NOT U102 ( .A(n118), .Z(n117) );
  GTECH_MUX2 U103 ( .A(n119), .B(n120), .S(n111), .Z(n118) );
  GTECH_NOT U104 ( .A(Mcand[2]), .Z(n111) );
  GTECH_NAND2 U105 ( .A(n121), .B(n86), .Z(n116) );
  GTECH_MUX2 U106 ( .A(n119), .B(n120), .S(Mcand[2]), .Z(n121) );
  GTECH_AOI22 U107 ( .A(n115), .B(n108), .C(n122), .D(n109), .Z(n120) );
  GTECH_AOI22 U108 ( .A(n113), .B(n108), .C(n110), .D(n109), .Z(n119) );
  GTECH_NOT U109 ( .A(n122), .Z(n110) );
  GTECH_OA21 U110 ( .A(Mcand[1]), .B(n123), .C(n124), .Z(n122) );
  GTECH_AO21 U111 ( .A(n123), .B(Mcand[1]), .C(n125), .Z(n124) );
  GTECH_NOT U112 ( .A(n17), .Z(n125) );
  GTECH_NOT U113 ( .A(n115), .Z(n113) );
  GTECH_OA21 U114 ( .A(Mcand[1]), .B(n90), .C(n126), .Z(n115) );
  GTECH_AO21 U115 ( .A(n90), .B(Mcand[1]), .C(n17), .Z(n126) );
  GTECH_MUX2 U116 ( .A(n127), .B(n128), .S(n17), .Z(N44) );
  GTECH_NOT U117 ( .A(n129), .Z(n128) );
  GTECH_MUX2 U118 ( .A(n130), .B(n131), .S(Mcand[1]), .Z(n129) );
  GTECH_NAND2 U119 ( .A(n132), .B(n86), .Z(n127) );
  GTECH_OR_NOT U120 ( .A(n93), .B(n14), .Z(n86) );
  GTECH_NOR2 U121 ( .A(n97), .B(n96), .Z(n93) );
  GTECH_MUX2 U122 ( .A(n131), .B(n130), .S(Mcand[1]), .Z(n132) );
  GTECH_AOI22 U123 ( .A(n123), .B(n109), .C(n90), .D(n108), .Z(n130) );
  GTECH_NOT U124 ( .A(n105), .Z(n108) );
  GTECH_NOT U125 ( .A(n107), .Z(n109) );
  GTECH_OA22 U126 ( .A(n123), .B(n107), .C(n90), .D(n105), .Z(n131) );
  GTECH_OR_NOT U127 ( .A(n14), .B(n96), .Z(n105) );
  GTECH_AND_NOT U128 ( .A(Mcand[0]), .B(n92), .Z(n90) );
  GTECH_OR_NOT U129 ( .A(n14), .B(n97), .Z(n107) );
  GTECH_AND2 U130 ( .A(Mcand[0]), .B(n92), .Z(n123) );
  GTECH_NOT U131 ( .A(n16), .Z(n92) );
  GTECH_OR_NOT U132 ( .A(n96), .B(n133), .Z(N42) );
  GTECH_NAND3 U133 ( .A(n134), .B(n135), .C(n97), .Z(n133) );
  GTECH_OA21 U134 ( .A(n12), .B(n85), .C(n97), .Z(N41) );
  GTECH_OAI21 U135 ( .A(n94), .B(n95), .C(n136), .Z(N40) );
  GTECH_AOI21 U136 ( .A(n12), .B(n97), .C(n96), .Z(n136) );
  GTECH_NOR3 U137 ( .A(n134), .B(n13), .C(n135), .Z(n96) );
  GTECH_AOI21 U138 ( .A(n12), .B(n85), .C(n137), .Z(n97) );
  GTECH_NOT U139 ( .A(St), .Z(n95) );
  GTECH_NOT U140 ( .A(n88), .Z(n94) );
  GTECH_NOR3 U141 ( .A(n135), .B(n134), .C(n137), .Z(n88) );
  GTECH_NOT U142 ( .A(n85), .Z(n135) );
  GTECH_AND3 U143 ( .A(n134), .B(n137), .C(n85), .Z(Done) );
  GTECH_NOT U144 ( .A(n13), .Z(n137) );
  GTECH_NOT U145 ( .A(n12), .Z(n134) );
endmodule

