
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI22 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NOT U83 ( .A(n97), .Z(n96) );
  GTECH_AND2 U84 ( .A(n93), .B(n94), .Z(n95) );
  GTECH_XOR2 U85 ( .A(n90), .B(n98), .Z(n86) );
  GTECH_NOT U86 ( .A(n89), .Z(n98) );
  GTECH_OAI22 U87 ( .A(n99), .B(n100), .C(n101), .D(n102), .Z(n89) );
  GTECH_AND2 U88 ( .A(n99), .B(n100), .Z(n101) );
  GTECH_NOT U89 ( .A(n103), .Z(n99) );
  GTECH_OR_NOT U90 ( .A(n104), .B(I_b[7]), .Z(n90) );
  GTECH_NOT U91 ( .A(n105), .Z(n84) );
  GTECH_OR_NOT U92 ( .A(n106), .B(n107), .Z(n105) );
  GTECH_XOR2 U93 ( .A(n108), .B(n107), .Z(N153) );
  GTECH_NOT U94 ( .A(n109), .Z(n107) );
  GTECH_XOR3 U95 ( .A(n110), .B(n93), .C(n97), .Z(n109) );
  GTECH_XOR3 U96 ( .A(n111), .B(n112), .C(n103), .Z(n97) );
  GTECH_OAI22 U97 ( .A(n113), .B(n114), .C(n115), .D(n116), .Z(n103) );
  GTECH_AND2 U98 ( .A(n113), .B(n114), .Z(n115) );
  GTECH_NOT U99 ( .A(n117), .Z(n113) );
  GTECH_NOT U100 ( .A(n102), .Z(n112) );
  GTECH_OR_NOT U101 ( .A(n118), .B(I_b[7]), .Z(n102) );
  GTECH_NOT U102 ( .A(n100), .Z(n111) );
  GTECH_OR_NOT U103 ( .A(n119), .B(I_a[7]), .Z(n100) );
  GTECH_NOT U104 ( .A(I_b[6]), .Z(n119) );
  GTECH_ADD_ABC U105 ( .A(n120), .B(n121), .C(n122), .COUT(n93) );
  GTECH_NOT U106 ( .A(n123), .Z(n122) );
  GTECH_XOR2 U107 ( .A(n124), .B(n125), .Z(n121) );
  GTECH_AND2 U108 ( .A(I_a[7]), .B(I_b[5]), .Z(n125) );
  GTECH_NOT U109 ( .A(n94), .Z(n110) );
  GTECH_OR_NOT U110 ( .A(n124), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U111 ( .A(n106), .Z(n108) );
  GTECH_OR_NOT U112 ( .A(n126), .B(n127), .Z(n106) );
  GTECH_XOR2 U113 ( .A(n126), .B(n128), .Z(N152) );
  GTECH_NOT U114 ( .A(n127), .Z(n128) );
  GTECH_XOR4 U115 ( .A(n129), .B(n124), .C(n120), .D(n123), .Z(n127) );
  GTECH_XOR3 U116 ( .A(n130), .B(n131), .C(n117), .Z(n123) );
  GTECH_OAI22 U117 ( .A(n132), .B(n133), .C(n134), .D(n135), .Z(n117) );
  GTECH_AND2 U118 ( .A(n132), .B(n133), .Z(n134) );
  GTECH_NOT U119 ( .A(n136), .Z(n132) );
  GTECH_NOT U120 ( .A(n116), .Z(n131) );
  GTECH_OR_NOT U121 ( .A(n137), .B(I_b[7]), .Z(n116) );
  GTECH_NOT U122 ( .A(n114), .Z(n130) );
  GTECH_OR_NOT U123 ( .A(n118), .B(I_b[6]), .Z(n114) );
  GTECH_NOT U124 ( .A(I_a[6]), .Z(n118) );
  GTECH_ADD_ABC U125 ( .A(n138), .B(n139), .C(n140), .COUT(n120) );
  GTECH_NOT U126 ( .A(n141), .Z(n140) );
  GTECH_XOR3 U127 ( .A(n142), .B(n143), .C(n144), .Z(n139) );
  GTECH_NOT U128 ( .A(n145), .Z(n142) );
  GTECH_OA21 U129 ( .A(n144), .B(n145), .C(n146), .Z(n124) );
  GTECH_AO21 U130 ( .A(n144), .B(n145), .C(n147), .Z(n146) );
  GTECH_NOT U131 ( .A(n148), .Z(n144) );
  GTECH_AND2 U132 ( .A(I_b[5]), .B(I_a[7]), .Z(n129) );
  GTECH_ADD_ABC U133 ( .A(n149), .B(n150), .C(n151), .COUT(n126) );
  GTECH_NOT U134 ( .A(n152), .Z(n151) );
  GTECH_OA22 U135 ( .A(n153), .B(n104), .C(n154), .D(n155), .Z(n150) );
  GTECH_OA21 U136 ( .A(n156), .B(n157), .C(n158), .Z(n149) );
  GTECH_AO21 U137 ( .A(n156), .B(n157), .C(n159), .Z(n158) );
  GTECH_XOR3 U138 ( .A(n160), .B(n152), .C(n161), .Z(N151) );
  GTECH_OA21 U139 ( .A(n156), .B(n157), .C(n162), .Z(n161) );
  GTECH_AO21 U140 ( .A(n156), .B(n157), .C(n159), .Z(n162) );
  GTECH_XOR2 U141 ( .A(n163), .B(n138), .Z(n152) );
  GTECH_ADD_ABC U142 ( .A(n164), .B(n165), .C(n166), .COUT(n138) );
  GTECH_NOT U143 ( .A(n167), .Z(n166) );
  GTECH_XOR3 U144 ( .A(n168), .B(n169), .C(n170), .Z(n165) );
  GTECH_XOR4 U145 ( .A(n143), .B(n148), .C(n145), .D(n141), .Z(n163) );
  GTECH_XOR3 U146 ( .A(n171), .B(n172), .C(n136), .Z(n141) );
  GTECH_OAI22 U147 ( .A(n173), .B(n174), .C(n175), .D(n176), .Z(n136) );
  GTECH_AND2 U148 ( .A(n173), .B(n174), .Z(n175) );
  GTECH_NOT U149 ( .A(n177), .Z(n173) );
  GTECH_NOT U150 ( .A(n135), .Z(n172) );
  GTECH_OR_NOT U151 ( .A(n178), .B(I_b[7]), .Z(n135) );
  GTECH_NOT U152 ( .A(n133), .Z(n171) );
  GTECH_OR_NOT U153 ( .A(n137), .B(I_b[6]), .Z(n133) );
  GTECH_NOT U154 ( .A(I_a[5]), .Z(n137) );
  GTECH_OR_NOT U155 ( .A(n179), .B(I_a[7]), .Z(n145) );
  GTECH_OAI22 U156 ( .A(n170), .B(n180), .C(n181), .D(n182), .Z(n148) );
  GTECH_AND2 U157 ( .A(n170), .B(n180), .Z(n181) );
  GTECH_NOT U158 ( .A(n183), .Z(n170) );
  GTECH_NOT U159 ( .A(n147), .Z(n143) );
  GTECH_OR_NOT U160 ( .A(n184), .B(I_a[6]), .Z(n147) );
  GTECH_OA22 U161 ( .A(n153), .B(n104), .C(n154), .D(n155), .Z(n160) );
  GTECH_NOT U162 ( .A(n185), .Z(n155) );
  GTECH_NOT U163 ( .A(I_a[7]), .Z(n104) );
  GTECH_XOR3 U164 ( .A(n156), .B(n186), .C(n159), .Z(N150) );
  GTECH_XOR2 U165 ( .A(n164), .B(n187), .Z(n159) );
  GTECH_XOR4 U166 ( .A(n169), .B(n183), .C(n167), .D(n168), .Z(n187) );
  GTECH_NOT U167 ( .A(n180), .Z(n168) );
  GTECH_OR_NOT U168 ( .A(n179), .B(I_a[6]), .Z(n180) );
  GTECH_XOR3 U169 ( .A(n188), .B(n189), .C(n177), .Z(n167) );
  GTECH_OAI22 U170 ( .A(n190), .B(n191), .C(n192), .D(n193), .Z(n177) );
  GTECH_AND2 U171 ( .A(n190), .B(n191), .Z(n192) );
  GTECH_NOT U172 ( .A(n194), .Z(n190) );
  GTECH_NOT U173 ( .A(n176), .Z(n189) );
  GTECH_OR_NOT U174 ( .A(n195), .B(I_b[7]), .Z(n176) );
  GTECH_NOT U175 ( .A(n174), .Z(n188) );
  GTECH_OR_NOT U176 ( .A(n178), .B(I_b[6]), .Z(n174) );
  GTECH_OAI22 U177 ( .A(n196), .B(n197), .C(n198), .D(n199), .Z(n183) );
  GTECH_AND2 U178 ( .A(n196), .B(n197), .Z(n198) );
  GTECH_NOT U179 ( .A(n182), .Z(n169) );
  GTECH_OR_NOT U180 ( .A(n184), .B(I_a[5]), .Z(n182) );
  GTECH_NOT U181 ( .A(I_b[5]), .Z(n184) );
  GTECH_ADD_ABC U182 ( .A(n200), .B(n201), .C(n202), .COUT(n164) );
  GTECH_NOT U183 ( .A(n203), .Z(n202) );
  GTECH_XOR3 U184 ( .A(n204), .B(n205), .C(n196), .Z(n201) );
  GTECH_NOT U185 ( .A(n206), .Z(n196) );
  GTECH_NOT U186 ( .A(n157), .Z(n186) );
  GTECH_XOR2 U187 ( .A(n185), .B(n154), .Z(n157) );
  GTECH_OA21 U188 ( .A(n207), .B(n208), .C(n209), .Z(n154) );
  GTECH_OR_NOT U189 ( .A(n210), .B(n211), .Z(n209) );
  GTECH_AND2 U190 ( .A(n207), .B(n208), .Z(n210) );
  GTECH_XOR2 U191 ( .A(n212), .B(n153), .Z(n185) );
  GTECH_OA21 U192 ( .A(n213), .B(n214), .C(n215), .Z(n153) );
  GTECH_AO21 U193 ( .A(n213), .B(n214), .C(n216), .Z(n215) );
  GTECH_NOT U194 ( .A(n217), .Z(n213) );
  GTECH_OR_NOT U195 ( .A(n218), .B(I_a[7]), .Z(n212) );
  GTECH_OA21 U196 ( .A(n219), .B(n220), .C(n221), .Z(n156) );
  GTECH_AO21 U197 ( .A(n219), .B(n220), .C(n222), .Z(n221) );
  GTECH_XOR3 U198 ( .A(n219), .B(n223), .C(n222), .Z(N149) );
  GTECH_XOR2 U199 ( .A(n200), .B(n224), .Z(n222) );
  GTECH_XOR4 U200 ( .A(n205), .B(n206), .C(n203), .D(n204), .Z(n224) );
  GTECH_NOT U201 ( .A(n197), .Z(n204) );
  GTECH_OR_NOT U202 ( .A(n179), .B(I_a[5]), .Z(n197) );
  GTECH_NOT U203 ( .A(I_b[4]), .Z(n179) );
  GTECH_XOR3 U204 ( .A(n225), .B(n226), .C(n194), .Z(n203) );
  GTECH_AO21 U205 ( .A(n227), .B(n228), .C(n229), .Z(n194) );
  GTECH_NOT U206 ( .A(n230), .Z(n229) );
  GTECH_NOT U207 ( .A(n193), .Z(n226) );
  GTECH_OR_NOT U208 ( .A(n231), .B(I_b[7]), .Z(n193) );
  GTECH_NOT U209 ( .A(n191), .Z(n225) );
  GTECH_OR_NOT U210 ( .A(n195), .B(I_b[6]), .Z(n191) );
  GTECH_OAI22 U211 ( .A(n232), .B(n233), .C(n234), .D(n235), .Z(n206) );
  GTECH_AND2 U212 ( .A(n232), .B(n233), .Z(n234) );
  GTECH_NOT U213 ( .A(n199), .Z(n205) );
  GTECH_OR_NOT U214 ( .A(n178), .B(I_b[5]), .Z(n199) );
  GTECH_ADD_ABC U215 ( .A(n236), .B(n237), .C(n238), .COUT(n200) );
  GTECH_XOR3 U216 ( .A(n239), .B(n240), .C(n232), .Z(n237) );
  GTECH_NOT U217 ( .A(n241), .Z(n232) );
  GTECH_NOT U218 ( .A(n233), .Z(n239) );
  GTECH_OA21 U219 ( .A(n242), .B(n243), .C(n244), .Z(n236) );
  GTECH_AO21 U220 ( .A(n242), .B(n243), .C(n245), .Z(n244) );
  GTECH_NOT U221 ( .A(n220), .Z(n223) );
  GTECH_XOR3 U222 ( .A(n246), .B(n207), .C(n211), .Z(n220) );
  GTECH_XOR3 U223 ( .A(n247), .B(n248), .C(n217), .Z(n211) );
  GTECH_OAI22 U224 ( .A(n249), .B(n250), .C(n251), .D(n252), .Z(n217) );
  GTECH_AND2 U225 ( .A(n249), .B(n250), .Z(n251) );
  GTECH_NOT U226 ( .A(n253), .Z(n249) );
  GTECH_NOT U227 ( .A(n216), .Z(n248) );
  GTECH_OR_NOT U228 ( .A(n218), .B(I_a[6]), .Z(n216) );
  GTECH_NOT U229 ( .A(n214), .Z(n247) );
  GTECH_OR_NOT U230 ( .A(n254), .B(I_a[7]), .Z(n214) );
  GTECH_ADD_ABC U231 ( .A(n255), .B(n256), .C(n257), .COUT(n207) );
  GTECH_XOR2 U232 ( .A(n258), .B(n259), .Z(n256) );
  GTECH_AND2 U233 ( .A(I_a[7]), .B(I_b[1]), .Z(n259) );
  GTECH_NOT U234 ( .A(n208), .Z(n246) );
  GTECH_OR_NOT U235 ( .A(n258), .B(I_a[7]), .Z(n208) );
  GTECH_ADD_ABC U236 ( .A(n260), .B(n261), .C(n262), .COUT(n219) );
  GTECH_XOR3 U237 ( .A(n255), .B(n263), .C(n257), .Z(n261) );
  GTECH_NOT U238 ( .A(n264), .Z(n257) );
  GTECH_XOR2 U239 ( .A(n260), .B(n265), .Z(N148) );
  GTECH_XOR4 U240 ( .A(n263), .B(n264), .C(n262), .D(n255), .Z(n265) );
  GTECH_ADD_ABC U241 ( .A(n266), .B(n267), .C(n268), .COUT(n255) );
  GTECH_XOR3 U242 ( .A(n269), .B(n270), .C(n271), .Z(n267) );
  GTECH_XOR2 U243 ( .A(n272), .B(n273), .Z(n262) );
  GTECH_OA21 U244 ( .A(n242), .B(n243), .C(n274), .Z(n273) );
  GTECH_AO21 U245 ( .A(n242), .B(n243), .C(n245), .Z(n274) );
  GTECH_XOR4 U246 ( .A(n240), .B(n241), .C(n233), .D(n238), .Z(n272) );
  GTECH_XOR3 U247 ( .A(n228), .B(n227), .C(n230), .Z(n238) );
  GTECH_NAND3 U248 ( .A(I_b[6]), .B(I_a[1]), .C(n275), .Z(n230) );
  GTECH_NOT U249 ( .A(n276), .Z(n227) );
  GTECH_OR_NOT U250 ( .A(n277), .B(I_b[7]), .Z(n276) );
  GTECH_NOT U251 ( .A(n278), .Z(n228) );
  GTECH_OR_NOT U252 ( .A(n231), .B(I_b[6]), .Z(n278) );
  GTECH_OR_NOT U253 ( .A(n178), .B(I_b[4]), .Z(n233) );
  GTECH_OAI22 U254 ( .A(n279), .B(n280), .C(n281), .D(n282), .Z(n241) );
  GTECH_AND2 U255 ( .A(n279), .B(n280), .Z(n281) );
  GTECH_NOT U256 ( .A(n283), .Z(n279) );
  GTECH_NOT U257 ( .A(n235), .Z(n240) );
  GTECH_OR_NOT U258 ( .A(n195), .B(I_b[5]), .Z(n235) );
  GTECH_XOR3 U259 ( .A(n284), .B(n285), .C(n253), .Z(n264) );
  GTECH_OAI22 U260 ( .A(n286), .B(n287), .C(n288), .D(n289), .Z(n253) );
  GTECH_AND2 U261 ( .A(n286), .B(n287), .Z(n288) );
  GTECH_NOT U262 ( .A(n290), .Z(n286) );
  GTECH_NOT U263 ( .A(n252), .Z(n285) );
  GTECH_OR_NOT U264 ( .A(n218), .B(I_a[5]), .Z(n252) );
  GTECH_NOT U265 ( .A(I_b[3]), .Z(n218) );
  GTECH_NOT U266 ( .A(n250), .Z(n284) );
  GTECH_OR_NOT U267 ( .A(n254), .B(I_a[6]), .Z(n250) );
  GTECH_XOR2 U268 ( .A(n291), .B(n258), .Z(n263) );
  GTECH_OA21 U269 ( .A(n271), .B(n292), .C(n293), .Z(n258) );
  GTECH_AO21 U270 ( .A(n271), .B(n292), .C(n294), .Z(n293) );
  GTECH_NOT U271 ( .A(n295), .Z(n271) );
  GTECH_AND2 U272 ( .A(I_b[1]), .B(I_a[7]), .Z(n291) );
  GTECH_ADD_ABC U273 ( .A(n296), .B(n297), .C(n298), .COUT(n260) );
  GTECH_NOT U274 ( .A(n299), .Z(n298) );
  GTECH_XOR3 U275 ( .A(n266), .B(n300), .C(n268), .Z(n297) );
  GTECH_NOT U276 ( .A(n301), .Z(n268) );
  GTECH_NOT U277 ( .A(n302), .Z(n300) );
  GTECH_XOR2 U278 ( .A(n303), .B(n296), .Z(N147) );
  GTECH_ADD_ABC U279 ( .A(n304), .B(n305), .C(n306), .COUT(n296) );
  GTECH_XOR3 U280 ( .A(n307), .B(n308), .C(n309), .Z(n305) );
  GTECH_OA21 U281 ( .A(n310), .B(n311), .C(n312), .Z(n304) );
  GTECH_AO21 U282 ( .A(n310), .B(n311), .C(n313), .Z(n312) );
  GTECH_XOR4 U283 ( .A(n301), .B(n266), .C(n302), .D(n299), .Z(n303) );
  GTECH_XOR3 U284 ( .A(n314), .B(n243), .C(n242), .Z(n299) );
  GTECH_XOR2 U285 ( .A(n315), .B(n275), .Z(n242) );
  GTECH_NOT U286 ( .A(n316), .Z(n275) );
  GTECH_OR_NOT U287 ( .A(n317), .B(I_b[7]), .Z(n316) );
  GTECH_OR_NOT U288 ( .A(n277), .B(I_b[6]), .Z(n315) );
  GTECH_NOT U289 ( .A(n318), .Z(n243) );
  GTECH_XOR3 U290 ( .A(n319), .B(n320), .C(n283), .Z(n318) );
  GTECH_AO21 U291 ( .A(n321), .B(n322), .C(n323), .Z(n283) );
  GTECH_NOT U292 ( .A(n324), .Z(n323) );
  GTECH_NOT U293 ( .A(n282), .Z(n320) );
  GTECH_OR_NOT U294 ( .A(n231), .B(I_b[5]), .Z(n282) );
  GTECH_NOT U295 ( .A(n280), .Z(n319) );
  GTECH_OR_NOT U296 ( .A(n195), .B(I_b[4]), .Z(n280) );
  GTECH_NOT U297 ( .A(n245), .Z(n314) );
  GTECH_NAND3 U298 ( .A(I_a[0]), .B(n325), .C(I_b[6]), .Z(n245) );
  GTECH_NOT U299 ( .A(n326), .Z(n325) );
  GTECH_XOR3 U300 ( .A(n269), .B(n270), .C(n295), .Z(n302) );
  GTECH_OAI22 U301 ( .A(n327), .B(n328), .C(n329), .D(n330), .Z(n295) );
  GTECH_AND2 U302 ( .A(n327), .B(n328), .Z(n329) );
  GTECH_NOT U303 ( .A(n294), .Z(n270) );
  GTECH_OR_NOT U304 ( .A(n331), .B(I_a[6]), .Z(n294) );
  GTECH_NOT U305 ( .A(n292), .Z(n269) );
  GTECH_OR_NOT U306 ( .A(n332), .B(I_a[7]), .Z(n292) );
  GTECH_ADD_ABC U307 ( .A(n307), .B(n333), .C(n309), .COUT(n266) );
  GTECH_NOT U308 ( .A(n334), .Z(n309) );
  GTECH_XOR3 U309 ( .A(n335), .B(n336), .C(n327), .Z(n333) );
  GTECH_NOT U310 ( .A(n337), .Z(n327) );
  GTECH_XOR3 U311 ( .A(n338), .B(n339), .C(n290), .Z(n301) );
  GTECH_OAI22 U312 ( .A(n340), .B(n341), .C(n342), .D(n343), .Z(n290) );
  GTECH_AND2 U313 ( .A(n340), .B(n341), .Z(n342) );
  GTECH_NOT U314 ( .A(n344), .Z(n340) );
  GTECH_NOT U315 ( .A(n289), .Z(n339) );
  GTECH_OR_NOT U316 ( .A(n178), .B(I_b[3]), .Z(n289) );
  GTECH_NOT U317 ( .A(n287), .Z(n338) );
  GTECH_OR_NOT U318 ( .A(n254), .B(I_a[5]), .Z(n287) );
  GTECH_NOT U319 ( .A(I_b[2]), .Z(n254) );
  GTECH_XOR2 U320 ( .A(n345), .B(n346), .Z(N146) );
  GTECH_XOR4 U321 ( .A(n308), .B(n334), .C(n306), .D(n307), .Z(n346) );
  GTECH_ADD_ABC U322 ( .A(n347), .B(n348), .C(n349), .COUT(n307) );
  GTECH_NOT U323 ( .A(n350), .Z(n349) );
  GTECH_XOR3 U324 ( .A(n351), .B(n352), .C(n353), .Z(n348) );
  GTECH_XOR2 U325 ( .A(n326), .B(n354), .Z(n306) );
  GTECH_AND2 U326 ( .A(I_b[6]), .B(I_a[0]), .Z(n354) );
  GTECH_XOR3 U327 ( .A(n322), .B(n321), .C(n324), .Z(n326) );
  GTECH_NAND3 U328 ( .A(I_b[4]), .B(I_a[1]), .C(n355), .Z(n324) );
  GTECH_NOT U329 ( .A(n356), .Z(n321) );
  GTECH_OR_NOT U330 ( .A(n277), .B(I_b[5]), .Z(n356) );
  GTECH_NOT U331 ( .A(n357), .Z(n322) );
  GTECH_OR_NOT U332 ( .A(n231), .B(I_b[4]), .Z(n357) );
  GTECH_XOR3 U333 ( .A(n358), .B(n359), .C(n344), .Z(n334) );
  GTECH_OAI22 U334 ( .A(n360), .B(n361), .C(n362), .D(n363), .Z(n344) );
  GTECH_AND2 U335 ( .A(n360), .B(n361), .Z(n362) );
  GTECH_NOT U336 ( .A(n364), .Z(n360) );
  GTECH_NOT U337 ( .A(n343), .Z(n359) );
  GTECH_OR_NOT U338 ( .A(n195), .B(I_b[3]), .Z(n343) );
  GTECH_NOT U339 ( .A(n341), .Z(n358) );
  GTECH_OR_NOT U340 ( .A(n178), .B(I_b[2]), .Z(n341) );
  GTECH_NOT U341 ( .A(I_a[4]), .Z(n178) );
  GTECH_NOT U342 ( .A(n365), .Z(n308) );
  GTECH_XOR3 U343 ( .A(n335), .B(n336), .C(n337), .Z(n365) );
  GTECH_OAI22 U344 ( .A(n353), .B(n366), .C(n367), .D(n368), .Z(n337) );
  GTECH_AND2 U345 ( .A(n353), .B(n366), .Z(n367) );
  GTECH_NOT U346 ( .A(n369), .Z(n353) );
  GTECH_NOT U347 ( .A(n330), .Z(n336) );
  GTECH_OR_NOT U348 ( .A(n331), .B(I_a[5]), .Z(n330) );
  GTECH_NOT U349 ( .A(n328), .Z(n335) );
  GTECH_OR_NOT U350 ( .A(n332), .B(I_a[6]), .Z(n328) );
  GTECH_OA21 U351 ( .A(n310), .B(n311), .C(n370), .Z(n345) );
  GTECH_AO21 U352 ( .A(n310), .B(n311), .C(n313), .Z(n370) );
  GTECH_XOR3 U353 ( .A(n371), .B(n311), .C(n310), .Z(N145) );
  GTECH_XOR2 U354 ( .A(n372), .B(n355), .Z(n310) );
  GTECH_NOT U355 ( .A(n373), .Z(n355) );
  GTECH_OR_NOT U356 ( .A(n317), .B(I_b[5]), .Z(n373) );
  GTECH_OR_NOT U357 ( .A(n277), .B(I_b[4]), .Z(n372) );
  GTECH_XOR2 U358 ( .A(n347), .B(n374), .Z(n311) );
  GTECH_XOR4 U359 ( .A(n352), .B(n369), .C(n350), .D(n351), .Z(n374) );
  GTECH_NOT U360 ( .A(n366), .Z(n351) );
  GTECH_OR_NOT U361 ( .A(n332), .B(I_a[5]), .Z(n366) );
  GTECH_XOR3 U362 ( .A(n375), .B(n376), .C(n364), .Z(n350) );
  GTECH_AO21 U363 ( .A(n377), .B(n378), .C(n379), .Z(n364) );
  GTECH_NOT U364 ( .A(n380), .Z(n379) );
  GTECH_NOT U365 ( .A(n363), .Z(n376) );
  GTECH_OR_NOT U366 ( .A(n231), .B(I_b[3]), .Z(n363) );
  GTECH_NOT U367 ( .A(n361), .Z(n375) );
  GTECH_OR_NOT U368 ( .A(n195), .B(I_b[2]), .Z(n361) );
  GTECH_OAI22 U369 ( .A(n381), .B(n382), .C(n383), .D(n384), .Z(n369) );
  GTECH_AND2 U370 ( .A(n381), .B(n382), .Z(n383) );
  GTECH_NOT U371 ( .A(n368), .Z(n352) );
  GTECH_OR_NOT U372 ( .A(n331), .B(I_a[4]), .Z(n368) );
  GTECH_ADD_ABC U373 ( .A(n385), .B(n386), .C(n387), .COUT(n347) );
  GTECH_XOR3 U374 ( .A(n388), .B(n389), .C(n381), .Z(n386) );
  GTECH_NOT U375 ( .A(n390), .Z(n381) );
  GTECH_OA21 U376 ( .A(n391), .B(n392), .C(n393), .Z(n385) );
  GTECH_AO21 U377 ( .A(n391), .B(n392), .C(n394), .Z(n393) );
  GTECH_NOT U378 ( .A(n313), .Z(n371) );
  GTECH_NAND3 U379 ( .A(I_a[0]), .B(n395), .C(I_b[4]), .Z(n313) );
  GTECH_XOR2 U380 ( .A(n396), .B(n395), .Z(N144) );
  GTECH_XOR2 U381 ( .A(n397), .B(n398), .Z(n395) );
  GTECH_XOR4 U382 ( .A(n389), .B(n390), .C(n387), .D(n388), .Z(n398) );
  GTECH_NOT U383 ( .A(n382), .Z(n388) );
  GTECH_OR_NOT U384 ( .A(n332), .B(I_a[4]), .Z(n382) );
  GTECH_NOT U385 ( .A(I_b[0]), .Z(n332) );
  GTECH_XOR3 U386 ( .A(n378), .B(n377), .C(n380), .Z(n387) );
  GTECH_NAND3 U387 ( .A(I_b[2]), .B(I_a[1]), .C(n399), .Z(n380) );
  GTECH_NOT U388 ( .A(n400), .Z(n377) );
  GTECH_OR_NOT U389 ( .A(n277), .B(I_b[3]), .Z(n400) );
  GTECH_NOT U390 ( .A(n401), .Z(n378) );
  GTECH_OR_NOT U391 ( .A(n231), .B(I_b[2]), .Z(n401) );
  GTECH_OAI22 U392 ( .A(n402), .B(n403), .C(n404), .D(n405), .Z(n390) );
  GTECH_AND2 U393 ( .A(n402), .B(n403), .Z(n404) );
  GTECH_NOT U394 ( .A(n406), .Z(n402) );
  GTECH_NOT U395 ( .A(n384), .Z(n389) );
  GTECH_OR_NOT U396 ( .A(n331), .B(I_a[3]), .Z(n384) );
  GTECH_OA21 U397 ( .A(n391), .B(n392), .C(n407), .Z(n397) );
  GTECH_AO21 U398 ( .A(n391), .B(n392), .C(n394), .Z(n407) );
  GTECH_AND2 U399 ( .A(I_b[4]), .B(I_a[0]), .Z(n396) );
  GTECH_XOR3 U400 ( .A(n408), .B(n392), .C(n391), .Z(N143) );
  GTECH_XOR2 U401 ( .A(n409), .B(n399), .Z(n391) );
  GTECH_NOT U402 ( .A(n410), .Z(n399) );
  GTECH_OR_NOT U403 ( .A(n317), .B(I_b[3]), .Z(n410) );
  GTECH_NOT U404 ( .A(I_a[0]), .Z(n317) );
  GTECH_OR_NOT U405 ( .A(n277), .B(I_b[2]), .Z(n409) );
  GTECH_NOT U406 ( .A(I_a[1]), .Z(n277) );
  GTECH_NOT U407 ( .A(n411), .Z(n392) );
  GTECH_XOR3 U408 ( .A(n412), .B(n413), .C(n406), .Z(n411) );
  GTECH_AO21 U409 ( .A(n414), .B(n415), .C(n416), .Z(n406) );
  GTECH_NOT U410 ( .A(n417), .Z(n416) );
  GTECH_NOT U411 ( .A(n405), .Z(n413) );
  GTECH_OR_NOT U412 ( .A(n231), .B(I_b[1]), .Z(n405) );
  GTECH_NOT U413 ( .A(n403), .Z(n412) );
  GTECH_OR_NOT U414 ( .A(n195), .B(I_b[0]), .Z(n403) );
  GTECH_NOT U415 ( .A(I_a[3]), .Z(n195) );
  GTECH_NOT U416 ( .A(n394), .Z(n408) );
  GTECH_NAND3 U417 ( .A(I_a[0]), .B(n418), .C(I_b[2]), .Z(n394) );
  GTECH_XOR2 U418 ( .A(n419), .B(n418), .Z(N142) );
  GTECH_NOT U419 ( .A(n420), .Z(n418) );
  GTECH_XOR3 U420 ( .A(n414), .B(n415), .C(n417), .Z(n420) );
  GTECH_NAND3 U421 ( .A(n421), .B(I_b[0]), .C(I_a[1]), .Z(n417) );
  GTECH_NOT U422 ( .A(n422), .Z(n415) );
  GTECH_OR_NOT U423 ( .A(n331), .B(I_a[1]), .Z(n422) );
  GTECH_NOT U424 ( .A(n423), .Z(n414) );
  GTECH_OR_NOT U425 ( .A(n231), .B(I_b[0]), .Z(n423) );
  GTECH_NOT U426 ( .A(I_a[2]), .Z(n231) );
  GTECH_AND2 U427 ( .A(I_b[2]), .B(I_a[0]), .Z(n419) );
  GTECH_XOR2 U428 ( .A(n421), .B(n424), .Z(N141) );
  GTECH_AND2 U429 ( .A(I_a[1]), .B(I_b[0]), .Z(n424) );
  GTECH_NOT U430 ( .A(n425), .Z(n421) );
  GTECH_OR_NOT U431 ( .A(n331), .B(I_a[0]), .Z(n425) );
  GTECH_NOT U432 ( .A(I_b[1]), .Z(n331) );
  GTECH_AND2 U433 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

