
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI21 U82 ( .A(n93), .B(n94), .C(n95), .Z(n87) );
  GTECH_OAI21 U83 ( .A(n96), .B(n97), .C(n98), .Z(n95) );
  GTECH_NOT U84 ( .A(n93), .Z(n97) );
  GTECH_XOR2 U85 ( .A(n90), .B(n99), .Z(n86) );
  GTECH_NOT U86 ( .A(n89), .Z(n99) );
  GTECH_OAI21 U87 ( .A(n100), .B(n101), .C(n102), .Z(n89) );
  GTECH_OAI21 U88 ( .A(n103), .B(n104), .C(n105), .Z(n102) );
  GTECH_NOT U89 ( .A(n104), .Z(n100) );
  GTECH_OR2 U90 ( .A(n106), .B(n107), .Z(n90) );
  GTECH_NOT U91 ( .A(n108), .Z(n84) );
  GTECH_OR2 U92 ( .A(n109), .B(n110), .Z(n108) );
  GTECH_XOR2 U93 ( .A(n111), .B(n112), .Z(N153) );
  GTECH_NOT U94 ( .A(n110), .Z(n112) );
  GTECH_XOR3 U95 ( .A(n96), .B(n93), .C(n98), .Z(n110) );
  GTECH_XOR3 U96 ( .A(n103), .B(n105), .C(n104), .Z(n98) );
  GTECH_OAI21 U97 ( .A(n113), .B(n114), .C(n115), .Z(n104) );
  GTECH_OAI21 U98 ( .A(n116), .B(n117), .C(n118), .Z(n115) );
  GTECH_NOT U99 ( .A(n117), .Z(n113) );
  GTECH_NOT U100 ( .A(n119), .Z(n105) );
  GTECH_OR2 U101 ( .A(n120), .B(n107), .Z(n119) );
  GTECH_NOT U102 ( .A(n101), .Z(n103) );
  GTECH_OR2 U103 ( .A(n121), .B(n106), .Z(n101) );
  GTECH_ADD_ABC U104 ( .A(n122), .B(n123), .C(n124), .COUT(n93) );
  GTECH_NOT U105 ( .A(n125), .Z(n124) );
  GTECH_XOR2 U106 ( .A(n126), .B(n127), .Z(n123) );
  GTECH_AND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n127) );
  GTECH_NOT U108 ( .A(n94), .Z(n96) );
  GTECH_OR2 U109 ( .A(n126), .B(n106), .Z(n94) );
  GTECH_NOT U110 ( .A(n109), .Z(n111) );
  GTECH_OR2 U111 ( .A(n128), .B(n129), .Z(n109) );
  GTECH_XOR2 U112 ( .A(n128), .B(n129), .Z(N152) );
  GTECH_XOR4 U113 ( .A(n126), .B(n125), .C(n130), .D(n122), .Z(n129) );
  GTECH_ADD_ABC U114 ( .A(n131), .B(n132), .C(n133), .COUT(n122) );
  GTECH_NOT U115 ( .A(n134), .Z(n133) );
  GTECH_XOR3 U116 ( .A(n135), .B(n136), .C(n137), .Z(n132) );
  GTECH_OR2 U117 ( .A(n106), .B(n138), .Z(n130) );
  GTECH_XOR3 U118 ( .A(n116), .B(n118), .C(n117), .Z(n125) );
  GTECH_OAI21 U119 ( .A(n139), .B(n140), .C(n141), .Z(n117) );
  GTECH_OAI21 U120 ( .A(n142), .B(n143), .C(n144), .Z(n141) );
  GTECH_NOT U121 ( .A(n143), .Z(n139) );
  GTECH_NOT U122 ( .A(n145), .Z(n118) );
  GTECH_OR2 U123 ( .A(n146), .B(n107), .Z(n145) );
  GTECH_NOT U124 ( .A(n114), .Z(n116) );
  GTECH_OR2 U125 ( .A(n120), .B(n121), .Z(n114) );
  GTECH_OA21 U126 ( .A(n137), .B(n147), .C(n148), .Z(n126) );
  GTECH_OAI21 U127 ( .A(n135), .B(n149), .C(n136), .Z(n148) );
  GTECH_NOT U128 ( .A(n147), .Z(n135) );
  GTECH_NOT U129 ( .A(n149), .Z(n137) );
  GTECH_ADD_ABC U130 ( .A(n150), .B(n151), .C(n152), .COUT(n128) );
  GTECH_NOT U131 ( .A(n153), .Z(n152) );
  GTECH_OA22 U132 ( .A(n154), .B(n106), .C(n155), .D(n156), .Z(n151) );
  GTECH_OA21 U133 ( .A(n157), .B(n158), .C(n159), .Z(n150) );
  GTECH_XOR3 U134 ( .A(n160), .B(n153), .C(n161), .Z(N151) );
  GTECH_OA21 U135 ( .A(n157), .B(n158), .C(n159), .Z(n161) );
  GTECH_OAI21 U136 ( .A(n162), .B(n163), .C(n164), .Z(n159) );
  GTECH_XOR2 U137 ( .A(n165), .B(n131), .Z(n153) );
  GTECH_ADD_ABC U138 ( .A(n166), .B(n167), .C(n168), .COUT(n131) );
  GTECH_NOT U139 ( .A(n169), .Z(n168) );
  GTECH_XOR3 U140 ( .A(n170), .B(n171), .C(n172), .Z(n167) );
  GTECH_XOR4 U141 ( .A(n136), .B(n149), .C(n147), .D(n134), .Z(n165) );
  GTECH_XOR3 U142 ( .A(n142), .B(n144), .C(n143), .Z(n134) );
  GTECH_OAI21 U143 ( .A(n173), .B(n174), .C(n175), .Z(n143) );
  GTECH_OAI21 U144 ( .A(n176), .B(n177), .C(n178), .Z(n175) );
  GTECH_NOT U145 ( .A(n177), .Z(n173) );
  GTECH_NOT U146 ( .A(n179), .Z(n144) );
  GTECH_OR2 U147 ( .A(n180), .B(n107), .Z(n179) );
  GTECH_NOT U148 ( .A(n140), .Z(n142) );
  GTECH_OR2 U149 ( .A(n146), .B(n121), .Z(n140) );
  GTECH_OR2 U150 ( .A(n181), .B(n106), .Z(n147) );
  GTECH_OAI21 U151 ( .A(n172), .B(n182), .C(n183), .Z(n149) );
  GTECH_OAI21 U152 ( .A(n170), .B(n184), .C(n171), .Z(n183) );
  GTECH_NOT U153 ( .A(n182), .Z(n170) );
  GTECH_NOT U154 ( .A(n184), .Z(n172) );
  GTECH_NOT U155 ( .A(n185), .Z(n136) );
  GTECH_OR2 U156 ( .A(n138), .B(n120), .Z(n185) );
  GTECH_OA22 U157 ( .A(n154), .B(n106), .C(n155), .D(n156), .Z(n160) );
  GTECH_NOT U158 ( .A(n186), .Z(n156) );
  GTECH_XOR3 U159 ( .A(n157), .B(n162), .C(n187), .Z(N150) );
  GTECH_NOT U160 ( .A(n164), .Z(n187) );
  GTECH_XOR2 U161 ( .A(n188), .B(n166), .Z(n164) );
  GTECH_ADD_ABC U162 ( .A(n189), .B(n190), .C(n191), .COUT(n166) );
  GTECH_NOT U163 ( .A(n192), .Z(n191) );
  GTECH_XOR3 U164 ( .A(n193), .B(n194), .C(n195), .Z(n190) );
  GTECH_XOR4 U165 ( .A(n171), .B(n184), .C(n182), .D(n169), .Z(n188) );
  GTECH_XOR3 U166 ( .A(n176), .B(n178), .C(n177), .Z(n169) );
  GTECH_OAI21 U167 ( .A(n196), .B(n197), .C(n198), .Z(n177) );
  GTECH_OAI21 U168 ( .A(n199), .B(n200), .C(n201), .Z(n198) );
  GTECH_NOT U169 ( .A(n200), .Z(n196) );
  GTECH_NOT U170 ( .A(n202), .Z(n178) );
  GTECH_OR2 U171 ( .A(n203), .B(n107), .Z(n202) );
  GTECH_NOT U172 ( .A(n174), .Z(n176) );
  GTECH_OR2 U173 ( .A(n180), .B(n121), .Z(n174) );
  GTECH_OR2 U174 ( .A(n181), .B(n120), .Z(n182) );
  GTECH_OAI21 U175 ( .A(n195), .B(n204), .C(n205), .Z(n184) );
  GTECH_OAI21 U176 ( .A(n193), .B(n206), .C(n194), .Z(n205) );
  GTECH_NOT U177 ( .A(n204), .Z(n193) );
  GTECH_NOT U178 ( .A(n206), .Z(n195) );
  GTECH_NOT U179 ( .A(n207), .Z(n171) );
  GTECH_OR2 U180 ( .A(n138), .B(n146), .Z(n207) );
  GTECH_NOT U181 ( .A(n158), .Z(n162) );
  GTECH_XOR2 U182 ( .A(n186), .B(n155), .Z(n158) );
  GTECH_OA21 U183 ( .A(n208), .B(n209), .C(n210), .Z(n155) );
  GTECH_OAI21 U184 ( .A(n211), .B(n212), .C(n213), .Z(n210) );
  GTECH_NOT U185 ( .A(n208), .Z(n212) );
  GTECH_XOR2 U186 ( .A(n214), .B(n154), .Z(n186) );
  GTECH_OA21 U187 ( .A(n215), .B(n216), .C(n217), .Z(n154) );
  GTECH_OAI21 U188 ( .A(n218), .B(n219), .C(n220), .Z(n217) );
  GTECH_NOT U189 ( .A(n219), .Z(n216) );
  GTECH_OR2 U190 ( .A(n221), .B(n106), .Z(n214) );
  GTECH_NOT U191 ( .A(n163), .Z(n157) );
  GTECH_OAI21 U192 ( .A(n222), .B(n223), .C(n224), .Z(n163) );
  GTECH_OAI21 U193 ( .A(n225), .B(n226), .C(n227), .Z(n224) );
  GTECH_NOT U194 ( .A(n222), .Z(n226) );
  GTECH_XOR3 U195 ( .A(n222), .B(n225), .C(n228), .Z(N149) );
  GTECH_NOT U196 ( .A(n227), .Z(n228) );
  GTECH_XOR2 U197 ( .A(n229), .B(n189), .Z(n227) );
  GTECH_ADD_ABC U198 ( .A(n230), .B(n231), .C(n232), .COUT(n189) );
  GTECH_XOR3 U199 ( .A(n233), .B(n234), .C(n235), .Z(n231) );
  GTECH_OA21 U200 ( .A(n236), .B(n237), .C(n238), .Z(n230) );
  GTECH_XOR4 U201 ( .A(n194), .B(n206), .C(n204), .D(n192), .Z(n229) );
  GTECH_XOR3 U202 ( .A(n199), .B(n201), .C(n200), .Z(n192) );
  GTECH_OAI21 U203 ( .A(n239), .B(n240), .C(n241), .Z(n200) );
  GTECH_NOT U204 ( .A(n242), .Z(n201) );
  GTECH_OR2 U205 ( .A(n243), .B(n107), .Z(n242) );
  GTECH_NOT U206 ( .A(n197), .Z(n199) );
  GTECH_OR2 U207 ( .A(n203), .B(n121), .Z(n197) );
  GTECH_OR2 U208 ( .A(n181), .B(n146), .Z(n204) );
  GTECH_OAI21 U209 ( .A(n235), .B(n244), .C(n245), .Z(n206) );
  GTECH_OAI21 U210 ( .A(n233), .B(n246), .C(n234), .Z(n245) );
  GTECH_NOT U211 ( .A(n244), .Z(n233) );
  GTECH_NOT U212 ( .A(n246), .Z(n235) );
  GTECH_NOT U213 ( .A(n247), .Z(n194) );
  GTECH_OR2 U214 ( .A(n180), .B(n138), .Z(n247) );
  GTECH_NOT U215 ( .A(n223), .Z(n225) );
  GTECH_XOR3 U216 ( .A(n211), .B(n208), .C(n213), .Z(n223) );
  GTECH_XOR3 U217 ( .A(n218), .B(n220), .C(n219), .Z(n213) );
  GTECH_OAI21 U218 ( .A(n248), .B(n249), .C(n250), .Z(n219) );
  GTECH_OAI21 U219 ( .A(n251), .B(n252), .C(n253), .Z(n250) );
  GTECH_NOT U220 ( .A(n252), .Z(n248) );
  GTECH_NOT U221 ( .A(n254), .Z(n220) );
  GTECH_OR2 U222 ( .A(n221), .B(n120), .Z(n254) );
  GTECH_NOT U223 ( .A(n215), .Z(n218) );
  GTECH_OR2 U224 ( .A(n255), .B(n106), .Z(n215) );
  GTECH_ADD_ABC U225 ( .A(n256), .B(n257), .C(n258), .COUT(n208) );
  GTECH_XOR2 U226 ( .A(n259), .B(n260), .Z(n257) );
  GTECH_AND2 U227 ( .A(I_a[7]), .B(I_b[1]), .Z(n260) );
  GTECH_NOT U228 ( .A(n209), .Z(n211) );
  GTECH_OR2 U229 ( .A(n259), .B(n106), .Z(n209) );
  GTECH_ADD_ABC U230 ( .A(n261), .B(n262), .C(n263), .COUT(n222) );
  GTECH_XOR3 U231 ( .A(n256), .B(n264), .C(n258), .Z(n262) );
  GTECH_NOT U232 ( .A(n265), .Z(n258) );
  GTECH_XOR2 U233 ( .A(n261), .B(n266), .Z(N148) );
  GTECH_XOR4 U234 ( .A(n264), .B(n265), .C(n263), .D(n256), .Z(n266) );
  GTECH_ADD_ABC U235 ( .A(n267), .B(n268), .C(n269), .COUT(n256) );
  GTECH_XOR3 U236 ( .A(n270), .B(n271), .C(n272), .Z(n268) );
  GTECH_XOR2 U237 ( .A(n273), .B(n274), .Z(n263) );
  GTECH_OA21 U238 ( .A(n236), .B(n237), .C(n238), .Z(n274) );
  GTECH_OAI21 U239 ( .A(n275), .B(n276), .C(n277), .Z(n238) );
  GTECH_NOT U240 ( .A(n236), .Z(n276) );
  GTECH_XOR4 U241 ( .A(n234), .B(n246), .C(n244), .D(n232), .Z(n273) );
  GTECH_XOR3 U242 ( .A(n278), .B(n279), .C(n241), .Z(n232) );
  GTECH_NAND3 U243 ( .A(I_b[7]), .B(I_a[0]), .C(n280), .Z(n241) );
  GTECH_NOT U244 ( .A(n240), .Z(n279) );
  GTECH_OR2 U245 ( .A(n281), .B(n107), .Z(n240) );
  GTECH_NOT U246 ( .A(n239), .Z(n278) );
  GTECH_OR2 U247 ( .A(n243), .B(n121), .Z(n239) );
  GTECH_OR2 U248 ( .A(n180), .B(n181), .Z(n244) );
  GTECH_OAI21 U249 ( .A(n282), .B(n283), .C(n284), .Z(n246) );
  GTECH_OAI21 U250 ( .A(n285), .B(n286), .C(n287), .Z(n284) );
  GTECH_NOT U251 ( .A(n286), .Z(n282) );
  GTECH_NOT U252 ( .A(n288), .Z(n234) );
  GTECH_OR2 U253 ( .A(n203), .B(n138), .Z(n288) );
  GTECH_XOR3 U254 ( .A(n251), .B(n253), .C(n252), .Z(n265) );
  GTECH_OAI21 U255 ( .A(n289), .B(n290), .C(n291), .Z(n252) );
  GTECH_OAI21 U256 ( .A(n292), .B(n293), .C(n294), .Z(n291) );
  GTECH_NOT U257 ( .A(n293), .Z(n289) );
  GTECH_NOT U258 ( .A(n295), .Z(n253) );
  GTECH_OR2 U259 ( .A(n221), .B(n146), .Z(n295) );
  GTECH_NOT U260 ( .A(n249), .Z(n251) );
  GTECH_OR2 U261 ( .A(n255), .B(n120), .Z(n249) );
  GTECH_XOR2 U262 ( .A(n296), .B(n259), .Z(n264) );
  GTECH_OA21 U263 ( .A(n272), .B(n297), .C(n298), .Z(n259) );
  GTECH_OAI21 U264 ( .A(n270), .B(n299), .C(n271), .Z(n298) );
  GTECH_NOT U265 ( .A(n299), .Z(n272) );
  GTECH_AND2 U266 ( .A(I_b[1]), .B(I_a[7]), .Z(n296) );
  GTECH_ADD_ABC U267 ( .A(n300), .B(n301), .C(n302), .COUT(n261) );
  GTECH_NOT U268 ( .A(n303), .Z(n302) );
  GTECH_XOR3 U269 ( .A(n267), .B(n304), .C(n269), .Z(n301) );
  GTECH_NOT U270 ( .A(n305), .Z(n269) );
  GTECH_NOT U271 ( .A(n306), .Z(n304) );
  GTECH_XOR2 U272 ( .A(n307), .B(n300), .Z(N147) );
  GTECH_ADD_ABC U273 ( .A(n308), .B(n309), .C(n310), .COUT(n300) );
  GTECH_XOR3 U274 ( .A(n311), .B(n312), .C(n313), .Z(n309) );
  GTECH_OA21 U275 ( .A(n314), .B(n315), .C(n316), .Z(n308) );
  GTECH_XOR4 U276 ( .A(n305), .B(n267), .C(n306), .D(n303), .Z(n307) );
  GTECH_XOR3 U277 ( .A(n277), .B(n237), .C(n236), .Z(n303) );
  GTECH_XOR2 U278 ( .A(n317), .B(n280), .Z(n236) );
  GTECH_NOT U279 ( .A(n318), .Z(n280) );
  GTECH_OR2 U280 ( .A(n281), .B(n121), .Z(n318) );
  GTECH_NOT U281 ( .A(I_b[6]), .Z(n121) );
  GTECH_OR2 U282 ( .A(n319), .B(n107), .Z(n317) );
  GTECH_NOT U283 ( .A(I_b[7]), .Z(n107) );
  GTECH_NOT U284 ( .A(n275), .Z(n237) );
  GTECH_XOR3 U285 ( .A(n285), .B(n287), .C(n286), .Z(n275) );
  GTECH_OAI21 U286 ( .A(n320), .B(n321), .C(n322), .Z(n286) );
  GTECH_NOT U287 ( .A(n323), .Z(n287) );
  GTECH_OR2 U288 ( .A(n243), .B(n138), .Z(n323) );
  GTECH_NOT U289 ( .A(n283), .Z(n285) );
  GTECH_OR2 U290 ( .A(n203), .B(n181), .Z(n283) );
  GTECH_NOT U291 ( .A(n324), .Z(n277) );
  GTECH_NAND3 U292 ( .A(I_a[0]), .B(n325), .C(I_b[6]), .Z(n324) );
  GTECH_NOT U293 ( .A(n326), .Z(n325) );
  GTECH_XOR3 U294 ( .A(n270), .B(n271), .C(n299), .Z(n306) );
  GTECH_OAI21 U295 ( .A(n327), .B(n328), .C(n329), .Z(n299) );
  GTECH_OAI21 U296 ( .A(n330), .B(n331), .C(n332), .Z(n329) );
  GTECH_NOT U297 ( .A(n333), .Z(n271) );
  GTECH_OR2 U298 ( .A(n334), .B(n120), .Z(n333) );
  GTECH_NOT U299 ( .A(n297), .Z(n270) );
  GTECH_OR2 U300 ( .A(n335), .B(n106), .Z(n297) );
  GTECH_NOT U301 ( .A(I_a[7]), .Z(n106) );
  GTECH_ADD_ABC U302 ( .A(n311), .B(n336), .C(n313), .COUT(n267) );
  GTECH_NOT U303 ( .A(n337), .Z(n313) );
  GTECH_XOR3 U304 ( .A(n330), .B(n332), .C(n327), .Z(n336) );
  GTECH_NOT U305 ( .A(n331), .Z(n327) );
  GTECH_XOR3 U306 ( .A(n292), .B(n294), .C(n293), .Z(n305) );
  GTECH_OAI21 U307 ( .A(n338), .B(n339), .C(n340), .Z(n293) );
  GTECH_OAI21 U308 ( .A(n341), .B(n342), .C(n343), .Z(n340) );
  GTECH_NOT U309 ( .A(n342), .Z(n338) );
  GTECH_NOT U310 ( .A(n344), .Z(n294) );
  GTECH_OR2 U311 ( .A(n180), .B(n221), .Z(n344) );
  GTECH_NOT U312 ( .A(n290), .Z(n292) );
  GTECH_OR2 U313 ( .A(n255), .B(n146), .Z(n290) );
  GTECH_XOR2 U314 ( .A(n345), .B(n346), .Z(N146) );
  GTECH_XOR4 U315 ( .A(n312), .B(n337), .C(n310), .D(n311), .Z(n346) );
  GTECH_ADD_ABC U316 ( .A(n347), .B(n348), .C(n349), .COUT(n311) );
  GTECH_NOT U317 ( .A(n350), .Z(n349) );
  GTECH_XOR3 U318 ( .A(n351), .B(n352), .C(n353), .Z(n348) );
  GTECH_XOR2 U319 ( .A(n326), .B(n354), .Z(n310) );
  GTECH_AND2 U320 ( .A(I_b[6]), .B(I_a[0]), .Z(n354) );
  GTECH_XOR3 U321 ( .A(n355), .B(n356), .C(n322), .Z(n326) );
  GTECH_NAND3 U322 ( .A(I_b[5]), .B(I_a[0]), .C(n357), .Z(n322) );
  GTECH_NOT U323 ( .A(n321), .Z(n356) );
  GTECH_OR2 U324 ( .A(n281), .B(n138), .Z(n321) );
  GTECH_NOT U325 ( .A(n320), .Z(n355) );
  GTECH_OR2 U326 ( .A(n243), .B(n181), .Z(n320) );
  GTECH_XOR3 U327 ( .A(n341), .B(n343), .C(n342), .Z(n337) );
  GTECH_OAI21 U328 ( .A(n358), .B(n359), .C(n360), .Z(n342) );
  GTECH_OAI21 U329 ( .A(n361), .B(n362), .C(n363), .Z(n360) );
  GTECH_NOT U330 ( .A(n362), .Z(n358) );
  GTECH_NOT U331 ( .A(n364), .Z(n343) );
  GTECH_OR2 U332 ( .A(n203), .B(n221), .Z(n364) );
  GTECH_NOT U333 ( .A(n339), .Z(n341) );
  GTECH_OR2 U334 ( .A(n180), .B(n255), .Z(n339) );
  GTECH_NOT U335 ( .A(n365), .Z(n312) );
  GTECH_XOR3 U336 ( .A(n330), .B(n332), .C(n331), .Z(n365) );
  GTECH_OAI21 U337 ( .A(n353), .B(n366), .C(n367), .Z(n331) );
  GTECH_OAI21 U338 ( .A(n351), .B(n368), .C(n352), .Z(n367) );
  GTECH_NOT U339 ( .A(n366), .Z(n351) );
  GTECH_NOT U340 ( .A(n368), .Z(n353) );
  GTECH_NOT U341 ( .A(n369), .Z(n332) );
  GTECH_OR2 U342 ( .A(n334), .B(n146), .Z(n369) );
  GTECH_NOT U343 ( .A(n328), .Z(n330) );
  GTECH_OR2 U344 ( .A(n335), .B(n120), .Z(n328) );
  GTECH_NOT U345 ( .A(I_a[6]), .Z(n120) );
  GTECH_OA21 U346 ( .A(n314), .B(n315), .C(n316), .Z(n345) );
  GTECH_OAI21 U347 ( .A(n370), .B(n371), .C(n372), .Z(n316) );
  GTECH_NOT U348 ( .A(n314), .Z(n371) );
  GTECH_XOR3 U349 ( .A(n372), .B(n315), .C(n314), .Z(N145) );
  GTECH_XOR2 U350 ( .A(n373), .B(n357), .Z(n314) );
  GTECH_NOT U351 ( .A(n374), .Z(n357) );
  GTECH_OR2 U352 ( .A(n281), .B(n181), .Z(n374) );
  GTECH_NOT U353 ( .A(I_b[4]), .Z(n181) );
  GTECH_OR2 U354 ( .A(n319), .B(n138), .Z(n373) );
  GTECH_NOT U355 ( .A(I_b[5]), .Z(n138) );
  GTECH_NOT U356 ( .A(n370), .Z(n315) );
  GTECH_XOR2 U357 ( .A(n375), .B(n347), .Z(n370) );
  GTECH_ADD_ABC U358 ( .A(n376), .B(n377), .C(n378), .COUT(n347) );
  GTECH_XOR3 U359 ( .A(n379), .B(n380), .C(n381), .Z(n377) );
  GTECH_OA21 U360 ( .A(n382), .B(n383), .C(n384), .Z(n376) );
  GTECH_XOR4 U361 ( .A(n352), .B(n368), .C(n366), .D(n350), .Z(n375) );
  GTECH_XOR3 U362 ( .A(n361), .B(n363), .C(n362), .Z(n350) );
  GTECH_OAI21 U363 ( .A(n385), .B(n386), .C(n387), .Z(n362) );
  GTECH_NOT U364 ( .A(n388), .Z(n363) );
  GTECH_OR2 U365 ( .A(n243), .B(n221), .Z(n388) );
  GTECH_NOT U366 ( .A(n359), .Z(n361) );
  GTECH_OR2 U367 ( .A(n203), .B(n255), .Z(n359) );
  GTECH_OR2 U368 ( .A(n335), .B(n146), .Z(n366) );
  GTECH_NOT U369 ( .A(I_a[5]), .Z(n146) );
  GTECH_OAI21 U370 ( .A(n381), .B(n389), .C(n390), .Z(n368) );
  GTECH_OAI21 U371 ( .A(n379), .B(n391), .C(n380), .Z(n390) );
  GTECH_NOT U372 ( .A(n391), .Z(n381) );
  GTECH_NOT U373 ( .A(n392), .Z(n352) );
  GTECH_OR2 U374 ( .A(n334), .B(n180), .Z(n392) );
  GTECH_NOT U375 ( .A(n393), .Z(n372) );
  GTECH_NAND3 U376 ( .A(I_a[0]), .B(n394), .C(I_b[4]), .Z(n393) );
  GTECH_XOR2 U377 ( .A(n395), .B(n394), .Z(N144) );
  GTECH_XOR2 U378 ( .A(n396), .B(n397), .Z(n394) );
  GTECH_XOR4 U379 ( .A(n380), .B(n391), .C(n378), .D(n379), .Z(n397) );
  GTECH_NOT U380 ( .A(n389), .Z(n379) );
  GTECH_OR2 U381 ( .A(n335), .B(n180), .Z(n389) );
  GTECH_NOT U382 ( .A(I_a[4]), .Z(n180) );
  GTECH_XOR3 U383 ( .A(n398), .B(n399), .C(n387), .Z(n378) );
  GTECH_NAND3 U384 ( .A(I_b[3]), .B(I_a[0]), .C(n400), .Z(n387) );
  GTECH_NOT U385 ( .A(n386), .Z(n399) );
  GTECH_OR2 U386 ( .A(n281), .B(n221), .Z(n386) );
  GTECH_NOT U387 ( .A(n385), .Z(n398) );
  GTECH_OR2 U388 ( .A(n243), .B(n255), .Z(n385) );
  GTECH_OAI21 U389 ( .A(n401), .B(n402), .C(n403), .Z(n391) );
  GTECH_OAI21 U390 ( .A(n404), .B(n405), .C(n406), .Z(n403) );
  GTECH_NOT U391 ( .A(n405), .Z(n401) );
  GTECH_NOT U392 ( .A(n407), .Z(n380) );
  GTECH_OR2 U393 ( .A(n334), .B(n203), .Z(n407) );
  GTECH_OA21 U394 ( .A(n382), .B(n383), .C(n384), .Z(n396) );
  GTECH_OAI21 U395 ( .A(n408), .B(n409), .C(n410), .Z(n384) );
  GTECH_NOT U396 ( .A(n382), .Z(n409) );
  GTECH_AND2 U397 ( .A(I_b[4]), .B(I_a[0]), .Z(n395) );
  GTECH_XOR3 U398 ( .A(n410), .B(n383), .C(n382), .Z(N143) );
  GTECH_XOR2 U399 ( .A(n411), .B(n400), .Z(n382) );
  GTECH_NOT U400 ( .A(n412), .Z(n400) );
  GTECH_OR2 U401 ( .A(n281), .B(n255), .Z(n412) );
  GTECH_NOT U402 ( .A(I_b[2]), .Z(n255) );
  GTECH_OR2 U403 ( .A(n319), .B(n221), .Z(n411) );
  GTECH_NOT U404 ( .A(I_b[3]), .Z(n221) );
  GTECH_NOT U405 ( .A(I_a[0]), .Z(n319) );
  GTECH_NOT U406 ( .A(n408), .Z(n383) );
  GTECH_XOR3 U407 ( .A(n404), .B(n406), .C(n405), .Z(n408) );
  GTECH_OAI21 U408 ( .A(n413), .B(n414), .C(n415), .Z(n405) );
  GTECH_NOT U409 ( .A(n416), .Z(n406) );
  GTECH_OR2 U410 ( .A(n243), .B(n334), .Z(n416) );
  GTECH_NOT U411 ( .A(n402), .Z(n404) );
  GTECH_OR2 U412 ( .A(n203), .B(n335), .Z(n402) );
  GTECH_NOT U413 ( .A(I_a[3]), .Z(n203) );
  GTECH_NOT U414 ( .A(n417), .Z(n410) );
  GTECH_NAND3 U415 ( .A(I_a[0]), .B(n418), .C(I_b[2]), .Z(n417) );
  GTECH_XOR2 U416 ( .A(n419), .B(n418), .Z(N142) );
  GTECH_NOT U417 ( .A(n420), .Z(n418) );
  GTECH_XOR3 U418 ( .A(n421), .B(n422), .C(n415), .Z(n420) );
  GTECH_NAND3 U419 ( .A(n423), .B(I_b[1]), .C(I_a[0]), .Z(n415) );
  GTECH_NOT U420 ( .A(n413), .Z(n422) );
  GTECH_OR2 U421 ( .A(n334), .B(n281), .Z(n413) );
  GTECH_NOT U422 ( .A(I_b[1]), .Z(n334) );
  GTECH_NOT U423 ( .A(n414), .Z(n421) );
  GTECH_OR2 U424 ( .A(n243), .B(n335), .Z(n414) );
  GTECH_NOT U425 ( .A(I_a[2]), .Z(n243) );
  GTECH_AND2 U426 ( .A(I_b[2]), .B(I_a[0]), .Z(n419) );
  GTECH_XOR2 U427 ( .A(n423), .B(n424), .Z(N141) );
  GTECH_AND2 U428 ( .A(I_a[0]), .B(I_b[1]), .Z(n424) );
  GTECH_NOT U429 ( .A(n425), .Z(n423) );
  GTECH_OR2 U430 ( .A(n335), .B(n281), .Z(n425) );
  GTECH_NOT U431 ( .A(I_a[1]), .Z(n281) );
  GTECH_NOT U432 ( .A(I_b[0]), .Z(n335) );
  GTECH_AND2 U433 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

