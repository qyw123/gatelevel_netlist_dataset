
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379;

  GTECH_MUX2 U133 ( .A(n272), .B(n273), .S(n274), .Z(sum[9]) );
  GTECH_XNOR2 U134 ( .A(n275), .B(n276), .Z(n273) );
  GTECH_XOR2 U135 ( .A(n276), .B(n277), .Z(n272) );
  GTECH_AOI21 U136 ( .A(a[9]), .B(b[9]), .C(n278), .Z(n276) );
  GTECH_NAND2 U137 ( .A(n279), .B(n280), .Z(sum[8]) );
  GTECH_OAI21 U138 ( .A(n281), .B(n282), .C(n283), .Z(n280) );
  GTECH_MUX2 U139 ( .A(n284), .B(n285), .S(n286), .Z(sum[7]) );
  GTECH_XOR2 U140 ( .A(n287), .B(n288), .Z(n285) );
  GTECH_OA21 U141 ( .A(a[6]), .B(n289), .C(n290), .Z(n287) );
  GTECH_AO21 U142 ( .A(n289), .B(a[6]), .C(b[6]), .Z(n290) );
  GTECH_XOR2 U143 ( .A(n288), .B(n291), .Z(n284) );
  GTECH_XOR2 U144 ( .A(a[7]), .B(b[7]), .Z(n288) );
  GTECH_MUX2 U145 ( .A(n292), .B(n293), .S(n294), .Z(sum[6]) );
  GTECH_XOR2 U146 ( .A(n295), .B(n296), .Z(n293) );
  GTECH_XNOR2 U147 ( .A(n295), .B(n289), .Z(n292) );
  GTECH_OAI21 U148 ( .A(n297), .B(n298), .C(n299), .Z(n289) );
  GTECH_XOR2 U149 ( .A(a[6]), .B(n300), .Z(n295) );
  GTECH_MUX2 U150 ( .A(n301), .B(n302), .S(n303), .Z(sum[5]) );
  GTECH_AND2 U151 ( .A(n304), .B(n299), .Z(n303) );
  GTECH_NOT U152 ( .A(n297), .Z(n304) );
  GTECH_AO21 U153 ( .A(n298), .B(n286), .C(n305), .Z(n302) );
  GTECH_OAI21 U154 ( .A(n305), .B(n286), .C(n298), .Z(n301) );
  GTECH_XOR2 U155 ( .A(n294), .B(n306), .Z(sum[4]) );
  GTECH_MUX2 U156 ( .A(n307), .B(n308), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U157 ( .A(n309), .B(n310), .Z(n308) );
  GTECH_XOR2 U158 ( .A(n311), .B(n309), .Z(n307) );
  GTECH_XOR2 U159 ( .A(a[3]), .B(b[3]), .Z(n309) );
  GTECH_OA21 U160 ( .A(a[2]), .B(n312), .C(n313), .Z(n311) );
  GTECH_AO21 U161 ( .A(n312), .B(a[2]), .C(b[2]), .Z(n313) );
  GTECH_MUX2 U162 ( .A(n314), .B(n315), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U163 ( .A(n316), .B(n317), .Z(n315) );
  GTECH_XNOR2 U164 ( .A(n316), .B(n312), .Z(n314) );
  GTECH_AO21 U165 ( .A(n318), .B(n319), .C(n320), .Z(n312) );
  GTECH_XOR2 U166 ( .A(a[2]), .B(n321), .Z(n316) );
  GTECH_MUX2 U167 ( .A(n322), .B(n323), .S(n324), .Z(sum[1]) );
  GTECH_AND2 U168 ( .A(n318), .B(n325), .Z(n324) );
  GTECH_OAI21 U169 ( .A(cin), .B(n319), .C(n326), .Z(n323) );
  GTECH_AO21 U170 ( .A(n326), .B(cin), .C(n319), .Z(n322) );
  GTECH_AND2 U171 ( .A(a[0]), .B(b[0]), .Z(n319) );
  GTECH_MUX2 U172 ( .A(n327), .B(n328), .S(n329), .Z(sum[15]) );
  GTECH_XOR2 U173 ( .A(n330), .B(n331), .Z(n328) );
  GTECH_ADD_ABC U174 ( .A(a[14]), .B(n332), .C(b[14]), .COUT(n330) );
  GTECH_XOR2 U175 ( .A(n331), .B(n333), .Z(n327) );
  GTECH_XOR2 U176 ( .A(a[15]), .B(b[15]), .Z(n331) );
  GTECH_MUX2 U177 ( .A(n334), .B(n335), .S(n329), .Z(sum[14]) );
  GTECH_XOR2 U178 ( .A(n332), .B(n336), .Z(n335) );
  GTECH_OA21 U179 ( .A(n337), .B(n338), .C(n339), .Z(n332) );
  GTECH_XOR2 U180 ( .A(n340), .B(n336), .Z(n334) );
  GTECH_XOR2 U181 ( .A(a[14]), .B(b[14]), .Z(n336) );
  GTECH_MUX2 U182 ( .A(n341), .B(n342), .S(n329), .Z(sum[13]) );
  GTECH_XOR2 U183 ( .A(n343), .B(n344), .Z(n342) );
  GTECH_XNOR2 U184 ( .A(n344), .B(n345), .Z(n341) );
  GTECH_OAI21 U185 ( .A(a[13]), .B(b[13]), .C(n346), .Z(n344) );
  GTECH_NOT U186 ( .A(n337), .Z(n346) );
  GTECH_NAND2 U187 ( .A(n347), .B(n348), .Z(sum[12]) );
  GTECH_OAI21 U188 ( .A(n338), .B(n349), .C(n350), .Z(n348) );
  GTECH_MUX2 U189 ( .A(n351), .B(n352), .S(n274), .Z(sum[11]) );
  GTECH_XOR2 U190 ( .A(n353), .B(n354), .Z(n352) );
  GTECH_AOI21 U191 ( .A(n355), .B(n356), .C(n357), .Z(n353) );
  GTECH_OA21 U192 ( .A(n356), .B(n355), .C(n358), .Z(n357) );
  GTECH_XOR2 U193 ( .A(n354), .B(n359), .Z(n351) );
  GTECH_XOR2 U194 ( .A(a[11]), .B(b[11]), .Z(n354) );
  GTECH_MUX2 U195 ( .A(n360), .B(n361), .S(n274), .Z(sum[10]) );
  GTECH_XOR2 U196 ( .A(n362), .B(n356), .Z(n361) );
  GTECH_AOI2N2 U197 ( .A(a[9]), .B(b[9]), .C(n278), .D(n275), .Z(n356) );
  GTECH_XOR2 U198 ( .A(n362), .B(n363), .Z(n360) );
  GTECH_XOR2 U199 ( .A(a[10]), .B(n358), .Z(n362) );
  GTECH_XOR2 U200 ( .A(cin), .B(n364), .Z(sum[0]) );
  GTECH_OAI21 U201 ( .A(n329), .B(n365), .C(n347), .Z(cout) );
  GTECH_NAND3 U202 ( .A(n343), .B(n345), .C(n329), .Z(n347) );
  GTECH_NOT U203 ( .A(n338), .Z(n343) );
  GTECH_AND2 U204 ( .A(b[12]), .B(a[12]), .Z(n338) );
  GTECH_AOI21 U205 ( .A(n333), .B(a[15]), .C(n366), .Z(n365) );
  GTECH_OA21 U206 ( .A(a[15]), .B(n333), .C(b[15]), .Z(n366) );
  GTECH_ADD_ABC U207 ( .A(a[14]), .B(n340), .C(b[14]), .COUT(n333) );
  GTECH_OA21 U208 ( .A(n337), .B(n345), .C(n339), .Z(n340) );
  GTECH_OR2 U209 ( .A(a[13]), .B(b[13]), .Z(n339) );
  GTECH_NOT U210 ( .A(n349), .Z(n345) );
  GTECH_NOR2 U211 ( .A(a[12]), .B(b[12]), .Z(n349) );
  GTECH_AND2 U212 ( .A(b[13]), .B(a[13]), .Z(n337) );
  GTECH_NOT U213 ( .A(n350), .Z(n329) );
  GTECH_OAI21 U214 ( .A(n367), .B(n274), .C(n279), .Z(n350) );
  GTECH_NAND3 U215 ( .A(n275), .B(n277), .C(n274), .Z(n279) );
  GTECH_NOT U216 ( .A(n281), .Z(n275) );
  GTECH_AND2 U217 ( .A(b[8]), .B(a[8]), .Z(n281) );
  GTECH_NOT U218 ( .A(n283), .Z(n274) );
  GTECH_MUX2 U219 ( .A(n368), .B(n306), .S(n286), .Z(n283) );
  GTECH_NOT U220 ( .A(n294), .Z(n286) );
  GTECH_MUX2 U221 ( .A(n364), .B(n369), .S(cin), .Z(n294) );
  GTECH_OA21 U222 ( .A(a[3]), .B(n310), .C(n370), .Z(n369) );
  GTECH_AO21 U223 ( .A(n310), .B(a[3]), .C(b[3]), .Z(n370) );
  GTECH_OAI21 U224 ( .A(n317), .B(n371), .C(n372), .Z(n310) );
  GTECH_AO21 U225 ( .A(n371), .B(n317), .C(n321), .Z(n372) );
  GTECH_NOT U226 ( .A(b[2]), .Z(n321) );
  GTECH_NOT U227 ( .A(a[2]), .Z(n371) );
  GTECH_AOI21 U228 ( .A(n318), .B(n326), .C(n320), .Z(n317) );
  GTECH_NOT U229 ( .A(n325), .Z(n320) );
  GTECH_NAND2 U230 ( .A(b[1]), .B(a[1]), .Z(n325) );
  GTECH_OR2 U231 ( .A(b[0]), .B(a[0]), .Z(n326) );
  GTECH_OR2 U232 ( .A(b[1]), .B(a[1]), .Z(n318) );
  GTECH_XOR2 U233 ( .A(a[0]), .B(b[0]), .Z(n364) );
  GTECH_AND2 U234 ( .A(n373), .B(n298), .Z(n306) );
  GTECH_NAND2 U235 ( .A(b[4]), .B(a[4]), .Z(n298) );
  GTECH_NOT U236 ( .A(n305), .Z(n373) );
  GTECH_OA21 U237 ( .A(a[7]), .B(n291), .C(n374), .Z(n368) );
  GTECH_AO21 U238 ( .A(n291), .B(a[7]), .C(b[7]), .Z(n374) );
  GTECH_OAI21 U239 ( .A(n296), .B(n375), .C(n376), .Z(n291) );
  GTECH_AO21 U240 ( .A(n375), .B(n296), .C(n300), .Z(n376) );
  GTECH_NOT U241 ( .A(b[6]), .Z(n300) );
  GTECH_NOT U242 ( .A(a[6]), .Z(n375) );
  GTECH_OA21 U243 ( .A(n305), .B(n297), .C(n299), .Z(n296) );
  GTECH_NAND2 U244 ( .A(b[5]), .B(a[5]), .Z(n299) );
  GTECH_NOR2 U245 ( .A(b[5]), .B(a[5]), .Z(n297) );
  GTECH_NOR2 U246 ( .A(b[4]), .B(a[4]), .Z(n305) );
  GTECH_AOI21 U247 ( .A(n359), .B(a[11]), .C(n377), .Z(n367) );
  GTECH_OA21 U248 ( .A(a[11]), .B(n359), .C(b[11]), .Z(n377) );
  GTECH_OAI21 U249 ( .A(n363), .B(n355), .C(n378), .Z(n359) );
  GTECH_AO21 U250 ( .A(n355), .B(n363), .C(n358), .Z(n378) );
  GTECH_NOT U251 ( .A(b[10]), .Z(n358) );
  GTECH_NOT U252 ( .A(a[10]), .Z(n355) );
  GTECH_AOI22 U253 ( .A(a[9]), .B(b[9]), .C(n277), .D(n379), .Z(n363) );
  GTECH_NOT U254 ( .A(n278), .Z(n379) );
  GTECH_NOR2 U255 ( .A(a[9]), .B(b[9]), .Z(n278) );
  GTECH_NOT U256 ( .A(n282), .Z(n277) );
  GTECH_NOR2 U257 ( .A(a[8]), .B(b[8]), .Z(n282) );
endmodule

