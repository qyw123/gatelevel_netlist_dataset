
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n113, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n113), .K(n113), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n250) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n113), .K(n113), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n113), .K(n113), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n113), .K(n113), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n113), .K(n113), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n113), .K(n113), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]), .QN(n267) );
  GTECH_FJK1S A_reg_15_ ( .J(n113), .K(n113), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n266) );
  GTECH_FJK1S A_reg_14_ ( .J(n113), .K(n113), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n265) );
  GTECH_FJK1S A_reg_13_ ( .J(n113), .K(n113), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n264) );
  GTECH_FJK1S A_reg_12_ ( .J(n113), .K(n113), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n263) );
  GTECH_FJK1S A_reg_11_ ( .J(n113), .K(n113), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n262) );
  GTECH_FJK1S A_reg_10_ ( .J(n113), .K(n113), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n261) );
  GTECH_FJK1S A_reg_9_ ( .J(n113), .K(n113), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n260) );
  GTECH_FJK1S A_reg_8_ ( .J(n113), .K(n113), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n259) );
  GTECH_FJK1S A_reg_7_ ( .J(n113), .K(n113), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n258) );
  GTECH_FJK1S A_reg_6_ ( .J(n113), .K(n113), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n257) );
  GTECH_FJK1S A_reg_5_ ( .J(n113), .K(n113), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n256) );
  GTECH_FJK1S A_reg_4_ ( .J(n113), .K(n113), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n255) );
  GTECH_FJK1S A_reg_3_ ( .J(n113), .K(n113), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n254) );
  GTECH_FJK1S A_reg_2_ ( .J(n113), .K(n113), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n253) );
  GTECH_FJK1S A_reg_1_ ( .J(n113), .K(n113), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n252) );
  GTECH_FJK1S A_reg_0_ ( .J(n113), .K(n113), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n251) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n113), .K(n113), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n113), .K(n113), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n113), .K(n113), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n113), .K(n113), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n113), .K(n113), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n113), .K(n113), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n113), .K(n113), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n113), .K(n113), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n113), .K(n113), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n113), .K(n113), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n113), .K(n113), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n113), .K(n113), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n113), .K(n113), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n113), .K(n113), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n113), .K(n113), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n113), .K(n113), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n113), .K(n113), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n113), .K(n113), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n113), .K(n113), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n113), .K(n113), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n113), .K(n113), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n113), .K(n113), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n113), .K(n113), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n113), .K(n113), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n113), .K(n113), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n113), .K(n113), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n113), .K(n113), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n113), .K(n113), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n113), .K(n113), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n113), .K(n113), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n113), .K(n113), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n113), .K(n113), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n113), .K(n113), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n113), .K(n113), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n113), .K(n113), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n113), .K(n113), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n113), .K(n113), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n113), .K(n113), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n113), .K(n113), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n113), .K(n113), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n113), .K(n113), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n113), .K(n113), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n113), .K(n113), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n113), .K(n113), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n113), .K(n113), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n113), .K(n113), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n113), .K(n113), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n113), .K(n113), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n113), .K(n113), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n113), .K(n113), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n113), .K(n113), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n113), .K(n113), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n113), .K(n113), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n113), .K(n113), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n113), .K(n113), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n113), .K(n113), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n113), .K(n113), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n113), .K(n113), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n113), .K(n113), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n113), .K(n113), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n113), .K(n113), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n113), .K(n113), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n113), .K(n113), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n113), .K(n113), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n113), .K(n113), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n113), .K(n113), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U252 ( .Z(n113) );
  GTECH_NOT U253 ( .A(n268), .Z(N99) );
  GTECH_AOI222 U254 ( .A(n269), .B(n270), .C(n271), .D(n272), .E(n273), .F(
        n274), .Z(n268) );
  GTECH_NOT U255 ( .A(n275), .Z(N98) );
  GTECH_AOI222 U256 ( .A(n271), .B(n276), .C(n277), .D(n278), .E(R[15]), .F(
        n279), .Z(n275) );
  GTECH_NAND2 U257 ( .A(n280), .B(n281), .Z(n277) );
  GTECH_OAI2N2 U258 ( .A(n13), .B(n282), .C(R[14]), .D(n279), .Z(N97) );
  GTECH_OAI2N2 U259 ( .A(n14), .B(n282), .C(R[13]), .D(n279), .Z(N96) );
  GTECH_OAI2N2 U260 ( .A(n15), .B(n282), .C(R[12]), .D(n279), .Z(N95) );
  GTECH_OAI2N2 U261 ( .A(n16), .B(n282), .C(R[11]), .D(n279), .Z(N94) );
  GTECH_OAI2N2 U262 ( .A(n17), .B(n282), .C(R[10]), .D(n279), .Z(N93) );
  GTECH_OAI2N2 U263 ( .A(n18), .B(n282), .C(R[9]), .D(n279), .Z(N92) );
  GTECH_OAI2N2 U264 ( .A(n19), .B(n282), .C(R[8]), .D(n279), .Z(N91) );
  GTECH_OAI2N2 U265 ( .A(n20), .B(n282), .C(R[7]), .D(n279), .Z(N90) );
  GTECH_OAI2N2 U266 ( .A(n21), .B(n282), .C(R[6]), .D(n279), .Z(N89) );
  GTECH_OAI2N2 U267 ( .A(n22), .B(n282), .C(R[5]), .D(n279), .Z(N88) );
  GTECH_OAI2N2 U268 ( .A(n23), .B(n282), .C(R[4]), .D(n279), .Z(N87) );
  GTECH_OAI2N2 U269 ( .A(n24), .B(n282), .C(R[3]), .D(n279), .Z(N86) );
  GTECH_OAI2N2 U270 ( .A(n25), .B(n282), .C(R[2]), .D(n279), .Z(N85) );
  GTECH_OAI2N2 U271 ( .A(n26), .B(n282), .C(R[1]), .D(n279), .Z(N84) );
  GTECH_OAI2N2 U272 ( .A(n27), .B(n282), .C(R[0]), .D(n279), .Z(N83) );
  GTECH_AND2 U273 ( .A(M[15]), .B(n279), .Z(N42) );
  GTECH_AND2 U274 ( .A(M[14]), .B(n279), .Z(N39) );
  GTECH_AND2 U275 ( .A(M[13]), .B(n279), .Z(N38) );
  GTECH_AND2 U276 ( .A(M[12]), .B(n279), .Z(N37) );
  GTECH_AND2 U277 ( .A(M[11]), .B(n279), .Z(N36) );
  GTECH_AND2 U278 ( .A(M[10]), .B(n279), .Z(N35) );
  GTECH_AND2 U279 ( .A(M[9]), .B(n279), .Z(N34) );
  GTECH_AND2 U280 ( .A(M[8]), .B(n279), .Z(N33) );
  GTECH_AND2 U281 ( .A(M[7]), .B(n279), .Z(N32) );
  GTECH_AND2 U282 ( .A(M[6]), .B(n279), .Z(N31) );
  GTECH_AND2 U283 ( .A(M[5]), .B(n279), .Z(N30) );
  GTECH_AND2 U284 ( .A(M[4]), .B(n279), .Z(N29) );
  GTECH_AND2 U285 ( .A(M[3]), .B(n279), .Z(N28) );
  GTECH_AND2 U286 ( .A(M[2]), .B(n279), .Z(N27) );
  GTECH_AND2 U287 ( .A(M[1]), .B(n279), .Z(N26) );
  GTECH_AND2 U288 ( .A(M[0]), .B(n279), .Z(N25) );
  GTECH_NOT U289 ( .A(n283), .Z(n279) );
  GTECH_NAND2 U290 ( .A(n283), .B(n284), .Z(N19) );
  GTECH_NAND3 U291 ( .A(n285), .B(n286), .C(n287), .Z(n284) );
  GTECH_NOT U292 ( .A(n9), .Z(n286) );
  GTECH_NAND3 U293 ( .A(n288), .B(n289), .C(n282), .Z(N18) );
  GTECH_OA21 U294 ( .A(n290), .B(n291), .C(n287), .Z(N17) );
  GTECH_AND_NOT U295 ( .A(n292), .B(n8), .Z(n290) );
  GTECH_OA21 U296 ( .A(n293), .B(n294), .C(n287), .Z(N16) );
  GTECH_AND_NOT U297 ( .A(n295), .B(n7), .Z(n293) );
  GTECH_NOT U298 ( .A(n296), .Z(N152) );
  GTECH_AOI222 U299 ( .A(n297), .B(n298), .C(n299), .D(n300), .E(n301), .F(
        n302), .Z(n296) );
  GTECH_NAND2 U300 ( .A(n289), .B(n303), .Z(N151) );
  GTECH_NOT U301 ( .A(n304), .Z(N150) );
  GTECH_AOI222 U302 ( .A(n305), .B(n297), .C(n299), .D(n306), .E(n301), .F(
        n307), .Z(n304) );
  GTECH_MUX2 U303 ( .A(n308), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND2 U304 ( .A(n287), .B(n309), .Z(n308) );
  GTECH_NOT U305 ( .A(n310), .Z(N149) );
  GTECH_AOI222 U306 ( .A(n311), .B(n297), .C(n299), .D(n312), .E(n301), .F(
        n313), .Z(n310) );
  GTECH_NOT U307 ( .A(n314), .Z(N148) );
  GTECH_AOI222 U308 ( .A(n315), .B(n297), .C(n299), .D(n316), .E(n301), .F(
        n317), .Z(n314) );
  GTECH_NOT U309 ( .A(n318), .Z(N147) );
  GTECH_AOI222 U310 ( .A(n319), .B(n297), .C(n299), .D(n320), .E(n301), .F(
        n321), .Z(n318) );
  GTECH_NOT U311 ( .A(n322), .Z(N146) );
  GTECH_AOI222 U312 ( .A(n323), .B(n297), .C(n299), .D(n324), .E(n301), .F(
        n325), .Z(n322) );
  GTECH_NOT U313 ( .A(n326), .Z(N145) );
  GTECH_AOI222 U314 ( .A(n327), .B(n297), .C(n299), .D(n328), .E(n301), .F(
        n329), .Z(n326) );
  GTECH_NOT U315 ( .A(n330), .Z(N144) );
  GTECH_AOI222 U316 ( .A(n331), .B(n297), .C(n299), .D(n332), .E(n301), .F(
        n333), .Z(n330) );
  GTECH_NOT U317 ( .A(n334), .Z(N143) );
  GTECH_AOI222 U318 ( .A(n335), .B(n297), .C(n299), .D(n336), .E(n301), .F(
        n337), .Z(n334) );
  GTECH_NOT U319 ( .A(n338), .Z(N142) );
  GTECH_AOI222 U320 ( .A(n339), .B(n297), .C(n299), .D(n340), .E(n301), .F(
        n341), .Z(n338) );
  GTECH_NOT U321 ( .A(n342), .Z(N141) );
  GTECH_AOI222 U322 ( .A(n343), .B(n297), .C(n299), .D(n344), .E(n301), .F(
        n345), .Z(n342) );
  GTECH_NOT U323 ( .A(n346), .Z(N140) );
  GTECH_AOI222 U324 ( .A(n347), .B(n297), .C(n299), .D(n348), .E(n301), .F(
        n349), .Z(n346) );
  GTECH_NOT U325 ( .A(n350), .Z(N14) );
  GTECH_NAND2 U326 ( .A(n287), .B(n250), .Z(n350) );
  GTECH_NOT U327 ( .A(n351), .Z(N139) );
  GTECH_AOI222 U328 ( .A(n352), .B(n297), .C(n299), .D(n353), .E(n301), .F(
        n354), .Z(n351) );
  GTECH_NOT U329 ( .A(n355), .Z(N138) );
  GTECH_AOI222 U330 ( .A(n356), .B(n297), .C(n299), .D(n357), .E(n301), .F(
        n358), .Z(n355) );
  GTECH_NOT U331 ( .A(n359), .Z(N137) );
  GTECH_AOI222 U332 ( .A(n360), .B(n297), .C(n299), .D(n361), .E(n301), .F(
        n362), .Z(n359) );
  GTECH_NOT U333 ( .A(n363), .Z(N136) );
  GTECH_AOI222 U334 ( .A(n297), .B(n270), .C(n299), .D(n272), .E(n301), .F(
        n274), .Z(n363) );
  GTECH_NOT U335 ( .A(n364), .Z(n274) );
  GTECH_XNOR2 U336 ( .A(n365), .B(n366), .Z(n364) );
  GTECH_NOT U337 ( .A(n367), .Z(n301) );
  GTECH_NOT U338 ( .A(n11), .Z(n272) );
  GTECH_NOT U339 ( .A(n368), .Z(n299) );
  GTECH_NOT U340 ( .A(n369), .Z(n270) );
  GTECH_XNOR2 U341 ( .A(n370), .B(n366), .Z(n369) );
  GTECH_NOT U342 ( .A(n371), .Z(n366) );
  GTECH_XNOR2 U343 ( .A(n252), .B(n11), .Z(n371) );
  GTECH_NOT U344 ( .A(n372), .Z(n370) );
  GTECH_NOT U345 ( .A(n373), .Z(n297) );
  GTECH_OAI2N2 U346 ( .A(n12), .B(n368), .C(n278), .D(n374), .Z(N135) );
  GTECH_NAND2 U347 ( .A(n373), .B(n367), .Z(n374) );
  GTECH_NAND3 U348 ( .A(n10), .B(n375), .C(N155), .Z(n367) );
  GTECH_NAND3 U349 ( .A(n28), .B(n376), .C(N155), .Z(n373) );
  GTECH_AO21 U350 ( .A(n251), .B(n276), .C(n365), .Z(n278) );
  GTECH_NAND2 U351 ( .A(n377), .B(N155), .Z(n368) );
  GTECH_XNOR2 U352 ( .A(n28), .B(n10), .Z(n377) );
  GTECH_AND2 U353 ( .A(N155), .B(n378), .Z(N134) );
  GTECH_NOT U354 ( .A(n13), .Z(n378) );
  GTECH_AND2 U355 ( .A(N155), .B(n379), .Z(N133) );
  GTECH_NOT U356 ( .A(n14), .Z(n379) );
  GTECH_AND2 U357 ( .A(N155), .B(n380), .Z(N132) );
  GTECH_NOT U358 ( .A(n15), .Z(n380) );
  GTECH_AND2 U359 ( .A(N155), .B(n381), .Z(N131) );
  GTECH_NOT U360 ( .A(n16), .Z(n381) );
  GTECH_AND2 U361 ( .A(N155), .B(n382), .Z(N130) );
  GTECH_NOT U362 ( .A(n17), .Z(n382) );
  GTECH_AND2 U363 ( .A(N155), .B(n383), .Z(N129) );
  GTECH_NOT U364 ( .A(n18), .Z(n383) );
  GTECH_AND2 U365 ( .A(N155), .B(n384), .Z(N128) );
  GTECH_NOT U366 ( .A(n19), .Z(n384) );
  GTECH_AND2 U367 ( .A(N155), .B(n385), .Z(N127) );
  GTECH_NOT U368 ( .A(n20), .Z(n385) );
  GTECH_AND2 U369 ( .A(N155), .B(n386), .Z(N126) );
  GTECH_NOT U370 ( .A(n21), .Z(n386) );
  GTECH_AND2 U371 ( .A(N155), .B(n387), .Z(N125) );
  GTECH_NOT U372 ( .A(n22), .Z(n387) );
  GTECH_AND2 U373 ( .A(N155), .B(n388), .Z(N124) );
  GTECH_NOT U374 ( .A(n23), .Z(n388) );
  GTECH_AND2 U375 ( .A(N155), .B(n389), .Z(N123) );
  GTECH_NOT U376 ( .A(n24), .Z(n389) );
  GTECH_AND2 U377 ( .A(N155), .B(n390), .Z(N122) );
  GTECH_NOT U378 ( .A(n25), .Z(n390) );
  GTECH_AND2 U379 ( .A(N155), .B(n391), .Z(N121) );
  GTECH_NOT U380 ( .A(n26), .Z(n391) );
  GTECH_AND2 U381 ( .A(N155), .B(n392), .Z(N120) );
  GTECH_NOT U382 ( .A(n27), .Z(n392) );
  GTECH_NOT U383 ( .A(n303), .Z(N155) );
  GTECH_NAND4 U384 ( .A(n8), .B(n7), .C(n9), .D(n393), .Z(n303) );
  GTECH_AND3 U385 ( .A(n289), .B(n309), .C(n6), .Z(n393) );
  GTECH_NOT U386 ( .A(n250), .Z(n309) );
  GTECH_NOT U387 ( .A(n394), .Z(N116) );
  GTECH_AOI222 U388 ( .A(n271), .B(n300), .C(n273), .D(n302), .E(n298), .F(
        n269), .Z(n394) );
  GTECH_XNOR2 U389 ( .A(n395), .B(n396), .Z(n298) );
  GTECH_NOT U390 ( .A(n397), .Z(n396) );
  GTECH_ADD_ABC U391 ( .A(n31), .B(n266), .C(n398), .COUT(n395) );
  GTECH_XNOR2 U392 ( .A(n399), .B(n397), .Z(n302) );
  GTECH_XNOR2 U393 ( .A(n30), .B(n267), .Z(n397) );
  GTECH_OA21 U394 ( .A(n400), .B(n31), .C(n401), .Z(n399) );
  GTECH_AO21 U395 ( .A(n31), .B(n400), .C(n402), .Z(n401) );
  GTECH_NOT U396 ( .A(n266), .Z(n400) );
  GTECH_NOT U397 ( .A(n30), .Z(n300) );
  GTECH_NAND2 U398 ( .A(n282), .B(n403), .Z(N115) );
  GTECH_NOT U399 ( .A(N41), .Z(n403) );
  GTECH_NAND2 U400 ( .A(n289), .B(n283), .Z(N41) );
  GTECH_NAND2 U401 ( .A(Ld), .B(n289), .Z(n283) );
  GTECH_NOT U402 ( .A(n404), .Z(N113) );
  GTECH_AOI222 U403 ( .A(n271), .B(n306), .C(n273), .D(n307), .E(n305), .F(
        n269), .Z(n404) );
  GTECH_XNOR2 U404 ( .A(n398), .B(n405), .Z(n305) );
  GTECH_ADD_ABC U405 ( .A(n32), .B(n265), .C(n406), .COUT(n398) );
  GTECH_NOT U406 ( .A(n407), .Z(n307) );
  GTECH_XNOR2 U407 ( .A(n402), .B(n405), .Z(n407) );
  GTECH_NOT U408 ( .A(n408), .Z(n405) );
  GTECH_XNOR2 U409 ( .A(n31), .B(n266), .Z(n408) );
  GTECH_OA21 U410 ( .A(n32), .B(n409), .C(n410), .Z(n402) );
  GTECH_AO21 U411 ( .A(n32), .B(n409), .C(n411), .Z(n410) );
  GTECH_NOT U412 ( .A(n265), .Z(n409) );
  GTECH_NOT U413 ( .A(n31), .Z(n306) );
  GTECH_NOT U414 ( .A(n412), .Z(N112) );
  GTECH_AOI222 U415 ( .A(n271), .B(n312), .C(n273), .D(n313), .E(n311), .F(
        n269), .Z(n412) );
  GTECH_XNOR2 U416 ( .A(n406), .B(n413), .Z(n311) );
  GTECH_ADD_ABC U417 ( .A(n33), .B(n264), .C(n414), .COUT(n406) );
  GTECH_NOT U418 ( .A(n415), .Z(n313) );
  GTECH_XNOR2 U419 ( .A(n411), .B(n413), .Z(n415) );
  GTECH_NOT U420 ( .A(n416), .Z(n413) );
  GTECH_XNOR2 U421 ( .A(n32), .B(n265), .Z(n416) );
  GTECH_OA21 U422 ( .A(n33), .B(n417), .C(n418), .Z(n411) );
  GTECH_AO21 U423 ( .A(n33), .B(n417), .C(n419), .Z(n418) );
  GTECH_NOT U424 ( .A(n264), .Z(n417) );
  GTECH_NOT U425 ( .A(n32), .Z(n312) );
  GTECH_NOT U426 ( .A(n420), .Z(N111) );
  GTECH_AOI222 U427 ( .A(n271), .B(n316), .C(n273), .D(n317), .E(n315), .F(
        n269), .Z(n420) );
  GTECH_XNOR2 U428 ( .A(n414), .B(n421), .Z(n315) );
  GTECH_ADD_ABC U429 ( .A(n34), .B(n263), .C(n422), .COUT(n414) );
  GTECH_NOT U430 ( .A(n423), .Z(n317) );
  GTECH_XNOR2 U431 ( .A(n419), .B(n421), .Z(n423) );
  GTECH_NOT U432 ( .A(n424), .Z(n421) );
  GTECH_XNOR2 U433 ( .A(n33), .B(n264), .Z(n424) );
  GTECH_OA21 U434 ( .A(n34), .B(n425), .C(n426), .Z(n419) );
  GTECH_AO21 U435 ( .A(n34), .B(n425), .C(n427), .Z(n426) );
  GTECH_NOT U436 ( .A(n263), .Z(n425) );
  GTECH_NOT U437 ( .A(n33), .Z(n316) );
  GTECH_NOT U438 ( .A(n428), .Z(N110) );
  GTECH_AOI222 U439 ( .A(n271), .B(n320), .C(n273), .D(n321), .E(n319), .F(
        n269), .Z(n428) );
  GTECH_XNOR2 U440 ( .A(n422), .B(n429), .Z(n319) );
  GTECH_ADD_ABC U441 ( .A(n35), .B(n262), .C(n430), .COUT(n422) );
  GTECH_NOT U442 ( .A(n431), .Z(n321) );
  GTECH_XNOR2 U443 ( .A(n427), .B(n429), .Z(n431) );
  GTECH_NOT U444 ( .A(n432), .Z(n429) );
  GTECH_XNOR2 U445 ( .A(n34), .B(n263), .Z(n432) );
  GTECH_OA21 U446 ( .A(n35), .B(n433), .C(n434), .Z(n427) );
  GTECH_AO21 U447 ( .A(n35), .B(n433), .C(n435), .Z(n434) );
  GTECH_NOT U448 ( .A(n262), .Z(n433) );
  GTECH_NOT U449 ( .A(n34), .Z(n320) );
  GTECH_NOT U450 ( .A(n436), .Z(N109) );
  GTECH_AOI222 U451 ( .A(n271), .B(n324), .C(n273), .D(n325), .E(n323), .F(
        n269), .Z(n436) );
  GTECH_XNOR2 U452 ( .A(n430), .B(n437), .Z(n323) );
  GTECH_ADD_ABC U453 ( .A(n36), .B(n261), .C(n438), .COUT(n430) );
  GTECH_NOT U454 ( .A(n439), .Z(n325) );
  GTECH_XNOR2 U455 ( .A(n435), .B(n437), .Z(n439) );
  GTECH_NOT U456 ( .A(n440), .Z(n437) );
  GTECH_XNOR2 U457 ( .A(n35), .B(n262), .Z(n440) );
  GTECH_OA21 U458 ( .A(n36), .B(n441), .C(n442), .Z(n435) );
  GTECH_AO21 U459 ( .A(n36), .B(n441), .C(n443), .Z(n442) );
  GTECH_NOT U460 ( .A(n261), .Z(n441) );
  GTECH_NOT U461 ( .A(n35), .Z(n324) );
  GTECH_NOT U462 ( .A(n444), .Z(N108) );
  GTECH_AOI222 U463 ( .A(n271), .B(n328), .C(n273), .D(n329), .E(n327), .F(
        n269), .Z(n444) );
  GTECH_XNOR2 U464 ( .A(n438), .B(n445), .Z(n327) );
  GTECH_ADD_ABC U465 ( .A(n37), .B(n260), .C(n446), .COUT(n438) );
  GTECH_NOT U466 ( .A(n447), .Z(n329) );
  GTECH_XNOR2 U467 ( .A(n443), .B(n445), .Z(n447) );
  GTECH_NOT U468 ( .A(n448), .Z(n445) );
  GTECH_XNOR2 U469 ( .A(n36), .B(n261), .Z(n448) );
  GTECH_OA21 U470 ( .A(n37), .B(n449), .C(n450), .Z(n443) );
  GTECH_AO21 U471 ( .A(n37), .B(n449), .C(n451), .Z(n450) );
  GTECH_NOT U472 ( .A(n260), .Z(n449) );
  GTECH_NOT U473 ( .A(n36), .Z(n328) );
  GTECH_NOT U474 ( .A(n452), .Z(N107) );
  GTECH_AOI222 U475 ( .A(n271), .B(n332), .C(n273), .D(n333), .E(n331), .F(
        n269), .Z(n452) );
  GTECH_XNOR2 U476 ( .A(n446), .B(n453), .Z(n331) );
  GTECH_ADD_ABC U477 ( .A(n38), .B(n259), .C(n454), .COUT(n446) );
  GTECH_NOT U478 ( .A(n455), .Z(n333) );
  GTECH_XNOR2 U479 ( .A(n451), .B(n453), .Z(n455) );
  GTECH_NOT U480 ( .A(n456), .Z(n453) );
  GTECH_XNOR2 U481 ( .A(n37), .B(n260), .Z(n456) );
  GTECH_OA21 U482 ( .A(n38), .B(n457), .C(n458), .Z(n451) );
  GTECH_AO21 U483 ( .A(n38), .B(n457), .C(n459), .Z(n458) );
  GTECH_NOT U484 ( .A(n259), .Z(n457) );
  GTECH_NOT U485 ( .A(n37), .Z(n332) );
  GTECH_NOT U486 ( .A(n460), .Z(N106) );
  GTECH_AOI222 U487 ( .A(n271), .B(n336), .C(n273), .D(n337), .E(n335), .F(
        n269), .Z(n460) );
  GTECH_XNOR2 U488 ( .A(n454), .B(n461), .Z(n335) );
  GTECH_ADD_ABC U489 ( .A(n39), .B(n258), .C(n462), .COUT(n454) );
  GTECH_NOT U490 ( .A(n463), .Z(n337) );
  GTECH_XNOR2 U491 ( .A(n459), .B(n461), .Z(n463) );
  GTECH_NOT U492 ( .A(n464), .Z(n461) );
  GTECH_XNOR2 U493 ( .A(n38), .B(n259), .Z(n464) );
  GTECH_OA21 U494 ( .A(n39), .B(n465), .C(n466), .Z(n459) );
  GTECH_AO21 U495 ( .A(n39), .B(n465), .C(n467), .Z(n466) );
  GTECH_NOT U496 ( .A(n258), .Z(n465) );
  GTECH_NOT U497 ( .A(n38), .Z(n336) );
  GTECH_NOT U498 ( .A(n468), .Z(N105) );
  GTECH_AOI222 U499 ( .A(n271), .B(n340), .C(n273), .D(n341), .E(n339), .F(
        n269), .Z(n468) );
  GTECH_XNOR2 U500 ( .A(n462), .B(n469), .Z(n339) );
  GTECH_ADD_ABC U501 ( .A(n40), .B(n257), .C(n470), .COUT(n462) );
  GTECH_NOT U502 ( .A(n471), .Z(n341) );
  GTECH_XNOR2 U503 ( .A(n467), .B(n469), .Z(n471) );
  GTECH_NOT U504 ( .A(n472), .Z(n469) );
  GTECH_XNOR2 U505 ( .A(n39), .B(n258), .Z(n472) );
  GTECH_OA21 U506 ( .A(n40), .B(n473), .C(n474), .Z(n467) );
  GTECH_AO21 U507 ( .A(n40), .B(n473), .C(n475), .Z(n474) );
  GTECH_NOT U508 ( .A(n257), .Z(n473) );
  GTECH_NOT U509 ( .A(n39), .Z(n340) );
  GTECH_NOT U510 ( .A(n476), .Z(N104) );
  GTECH_AOI222 U511 ( .A(n271), .B(n344), .C(n273), .D(n345), .E(n343), .F(
        n269), .Z(n476) );
  GTECH_XNOR2 U512 ( .A(n470), .B(n477), .Z(n343) );
  GTECH_ADD_ABC U513 ( .A(n41), .B(n256), .C(n478), .COUT(n470) );
  GTECH_NOT U514 ( .A(n479), .Z(n345) );
  GTECH_XNOR2 U515 ( .A(n475), .B(n477), .Z(n479) );
  GTECH_NOT U516 ( .A(n480), .Z(n477) );
  GTECH_XNOR2 U517 ( .A(n40), .B(n257), .Z(n480) );
  GTECH_OA21 U518 ( .A(n41), .B(n481), .C(n482), .Z(n475) );
  GTECH_AO21 U519 ( .A(n41), .B(n481), .C(n483), .Z(n482) );
  GTECH_NOT U520 ( .A(n256), .Z(n481) );
  GTECH_NOT U521 ( .A(n40), .Z(n344) );
  GTECH_NOT U522 ( .A(n484), .Z(N103) );
  GTECH_AOI222 U523 ( .A(n271), .B(n348), .C(n273), .D(n349), .E(n347), .F(
        n269), .Z(n484) );
  GTECH_XNOR2 U524 ( .A(n478), .B(n485), .Z(n347) );
  GTECH_ADD_ABC U525 ( .A(n42), .B(n255), .C(n486), .COUT(n478) );
  GTECH_NOT U526 ( .A(n487), .Z(n349) );
  GTECH_XNOR2 U527 ( .A(n483), .B(n485), .Z(n487) );
  GTECH_NOT U528 ( .A(n488), .Z(n485) );
  GTECH_XNOR2 U529 ( .A(n41), .B(n256), .Z(n488) );
  GTECH_OA21 U530 ( .A(n42), .B(n489), .C(n490), .Z(n483) );
  GTECH_AO21 U531 ( .A(n42), .B(n489), .C(n491), .Z(n490) );
  GTECH_NOT U532 ( .A(n255), .Z(n489) );
  GTECH_NOT U533 ( .A(n41), .Z(n348) );
  GTECH_NOT U534 ( .A(n492), .Z(N102) );
  GTECH_AOI222 U535 ( .A(n271), .B(n353), .C(n273), .D(n354), .E(n352), .F(
        n269), .Z(n492) );
  GTECH_XNOR2 U536 ( .A(n486), .B(n493), .Z(n352) );
  GTECH_ADD_ABC U537 ( .A(n43), .B(n254), .C(n494), .COUT(n486) );
  GTECH_NOT U538 ( .A(n495), .Z(n354) );
  GTECH_XNOR2 U539 ( .A(n491), .B(n493), .Z(n495) );
  GTECH_NOT U540 ( .A(n496), .Z(n493) );
  GTECH_XNOR2 U541 ( .A(n42), .B(n255), .Z(n496) );
  GTECH_OA21 U542 ( .A(n43), .B(n497), .C(n498), .Z(n491) );
  GTECH_AO21 U543 ( .A(n43), .B(n497), .C(n499), .Z(n498) );
  GTECH_NOT U544 ( .A(n254), .Z(n497) );
  GTECH_NOT U545 ( .A(n42), .Z(n353) );
  GTECH_NOT U546 ( .A(n500), .Z(N101) );
  GTECH_AOI222 U547 ( .A(n271), .B(n357), .C(n273), .D(n358), .E(n356), .F(
        n269), .Z(n500) );
  GTECH_XNOR2 U548 ( .A(n494), .B(n501), .Z(n356) );
  GTECH_ADD_ABC U549 ( .A(n29), .B(n253), .C(n502), .COUT(n494) );
  GTECH_NOT U550 ( .A(n503), .Z(n358) );
  GTECH_XNOR2 U551 ( .A(n499), .B(n501), .Z(n503) );
  GTECH_NOT U552 ( .A(n504), .Z(n501) );
  GTECH_XNOR2 U553 ( .A(n43), .B(n254), .Z(n504) );
  GTECH_OA21 U554 ( .A(n29), .B(n505), .C(n506), .Z(n499) );
  GTECH_AO21 U555 ( .A(n29), .B(n505), .C(n507), .Z(n506) );
  GTECH_NOT U556 ( .A(n253), .Z(n505) );
  GTECH_NOT U557 ( .A(n43), .Z(n357) );
  GTECH_NOT U558 ( .A(n508), .Z(N100) );
  GTECH_AOI222 U559 ( .A(n360), .B(n269), .C(n271), .D(n361), .E(n273), .F(
        n362), .Z(n508) );
  GTECH_NOT U560 ( .A(n509), .Z(n362) );
  GTECH_XNOR2 U561 ( .A(n507), .B(n510), .Z(n509) );
  GTECH_OA21 U562 ( .A(n11), .B(n511), .C(n512), .Z(n507) );
  GTECH_AO21 U563 ( .A(n11), .B(n511), .C(n365), .Z(n512) );
  GTECH_NOT U564 ( .A(n513), .Z(n365) );
  GTECH_NAND2 U565 ( .A(n12), .B(n514), .Z(n513) );
  GTECH_NOT U566 ( .A(n252), .Z(n511) );
  GTECH_NOT U567 ( .A(n281), .Z(n273) );
  GTECH_NAND2 U568 ( .A(N82), .B(n10), .Z(n281) );
  GTECH_NOT U569 ( .A(n515), .Z(N82) );
  GTECH_NOT U570 ( .A(n29), .Z(n361) );
  GTECH_NOT U571 ( .A(n516), .Z(n271) );
  GTECH_MUX2 U572 ( .A(n515), .B(n517), .S(n10), .Z(n516) );
  GTECH_NAND2 U573 ( .A(n28), .B(n287), .Z(n517) );
  GTECH_NAND2 U574 ( .A(n287), .B(n375), .Z(n515) );
  GTECH_NOT U575 ( .A(n28), .Z(n375) );
  GTECH_NOT U576 ( .A(n280), .Z(n269) );
  GTECH_NAND3 U577 ( .A(n287), .B(n376), .C(n28), .Z(n280) );
  GTECH_NOT U578 ( .A(n10), .Z(n376) );
  GTECH_NOT U579 ( .A(n282), .Z(n287) );
  GTECH_AO21 U580 ( .A(n9), .B(n291), .C(n518), .Z(n282) );
  GTECH_NAND2 U581 ( .A(n288), .B(n289), .Z(n518) );
  GTECH_NOT U582 ( .A(Rst), .Z(n289) );
  GTECH_NOT U583 ( .A(Ld), .Z(n288) );
  GTECH_NOT U584 ( .A(n285), .Z(n291) );
  GTECH_NAND2 U585 ( .A(n8), .B(n294), .Z(n285) );
  GTECH_NOT U586 ( .A(n292), .Z(n294) );
  GTECH_NAND2 U587 ( .A(n7), .B(n519), .Z(n292) );
  GTECH_NOT U588 ( .A(n295), .Z(n519) );
  GTECH_NAND2 U589 ( .A(n6), .B(n250), .Z(n295) );
  GTECH_XNOR2 U590 ( .A(n502), .B(n510), .Z(n360) );
  GTECH_NOT U591 ( .A(n520), .Z(n510) );
  GTECH_XNOR2 U592 ( .A(n29), .B(n253), .Z(n520) );
  GTECH_ADD_ABC U593 ( .A(n252), .B(n11), .C(n372), .COUT(n502) );
  GTECH_NAND2 U594 ( .A(n276), .B(n514), .Z(n372) );
  GTECH_NOT U595 ( .A(n251), .Z(n514) );
  GTECH_NOT U596 ( .A(n12), .Z(n276) );
endmodule

