
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI21 U82 ( .A(n93), .B(n94), .C(n95), .Z(n87) );
  GTECH_OAI21 U83 ( .A(n96), .B(n97), .C(n98), .Z(n95) );
  GTECH_NOT U84 ( .A(n93), .Z(n97) );
  GTECH_XOR2 U85 ( .A(n90), .B(n99), .Z(n86) );
  GTECH_NOT U86 ( .A(n89), .Z(n99) );
  GTECH_OAI21 U87 ( .A(n100), .B(n101), .C(n102), .Z(n89) );
  GTECH_OAI21 U88 ( .A(n103), .B(n104), .C(n105), .Z(n102) );
  GTECH_NOT U89 ( .A(n104), .Z(n100) );
  GTECH_OR_NOT U90 ( .A(n106), .B(I_b[7]), .Z(n90) );
  GTECH_NOT U91 ( .A(n107), .Z(n84) );
  GTECH_OR_NOT U92 ( .A(n108), .B(n109), .Z(n107) );
  GTECH_XOR2 U93 ( .A(n110), .B(n109), .Z(N153) );
  GTECH_NOT U94 ( .A(n111), .Z(n109) );
  GTECH_XOR3 U95 ( .A(n96), .B(n93), .C(n98), .Z(n111) );
  GTECH_XOR3 U96 ( .A(n103), .B(n105), .C(n104), .Z(n98) );
  GTECH_OAI21 U97 ( .A(n112), .B(n113), .C(n114), .Z(n104) );
  GTECH_OAI21 U98 ( .A(n115), .B(n116), .C(n117), .Z(n114) );
  GTECH_NOT U99 ( .A(n116), .Z(n112) );
  GTECH_NOT U100 ( .A(n118), .Z(n105) );
  GTECH_OR_NOT U101 ( .A(n119), .B(I_b[7]), .Z(n118) );
  GTECH_NOT U102 ( .A(n101), .Z(n103) );
  GTECH_OR_NOT U103 ( .A(n120), .B(I_a[7]), .Z(n101) );
  GTECH_NOT U104 ( .A(I_b[6]), .Z(n120) );
  GTECH_ADD_ABC U105 ( .A(n121), .B(n122), .C(n123), .COUT(n93) );
  GTECH_NOT U106 ( .A(n124), .Z(n123) );
  GTECH_XOR2 U107 ( .A(n125), .B(n126), .Z(n122) );
  GTECH_AND2 U108 ( .A(I_a[7]), .B(I_b[5]), .Z(n126) );
  GTECH_NOT U109 ( .A(n94), .Z(n96) );
  GTECH_OR_NOT U110 ( .A(n125), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U111 ( .A(n108), .Z(n110) );
  GTECH_OR_NOT U112 ( .A(n127), .B(n128), .Z(n108) );
  GTECH_XOR2 U113 ( .A(n127), .B(n129), .Z(N152) );
  GTECH_NOT U114 ( .A(n128), .Z(n129) );
  GTECH_XOR4 U115 ( .A(n130), .B(n125), .C(n121), .D(n124), .Z(n128) );
  GTECH_XOR3 U116 ( .A(n115), .B(n117), .C(n116), .Z(n124) );
  GTECH_OAI21 U117 ( .A(n131), .B(n132), .C(n133), .Z(n116) );
  GTECH_OAI21 U118 ( .A(n134), .B(n135), .C(n136), .Z(n133) );
  GTECH_NOT U119 ( .A(n135), .Z(n131) );
  GTECH_NOT U120 ( .A(n137), .Z(n117) );
  GTECH_OR_NOT U121 ( .A(n138), .B(I_b[7]), .Z(n137) );
  GTECH_NOT U122 ( .A(n113), .Z(n115) );
  GTECH_OR_NOT U123 ( .A(n119), .B(I_b[6]), .Z(n113) );
  GTECH_NOT U124 ( .A(I_a[6]), .Z(n119) );
  GTECH_ADD_ABC U125 ( .A(n139), .B(n140), .C(n141), .COUT(n121) );
  GTECH_NOT U126 ( .A(n142), .Z(n141) );
  GTECH_XOR3 U127 ( .A(n143), .B(n144), .C(n145), .Z(n140) );
  GTECH_OA21 U128 ( .A(n145), .B(n146), .C(n147), .Z(n125) );
  GTECH_OAI21 U129 ( .A(n143), .B(n148), .C(n144), .Z(n147) );
  GTECH_NOT U130 ( .A(n146), .Z(n143) );
  GTECH_NOT U131 ( .A(n148), .Z(n145) );
  GTECH_AND2 U132 ( .A(I_b[5]), .B(I_a[7]), .Z(n130) );
  GTECH_ADD_ABC U133 ( .A(n149), .B(n150), .C(n151), .COUT(n127) );
  GTECH_NOT U134 ( .A(n152), .Z(n151) );
  GTECH_OA22 U135 ( .A(n153), .B(n106), .C(n154), .D(n155), .Z(n150) );
  GTECH_OA21 U136 ( .A(n156), .B(n157), .C(n158), .Z(n149) );
  GTECH_XOR3 U137 ( .A(n159), .B(n152), .C(n160), .Z(N151) );
  GTECH_OA21 U138 ( .A(n156), .B(n157), .C(n158), .Z(n160) );
  GTECH_OAI21 U139 ( .A(n161), .B(n162), .C(n163), .Z(n158) );
  GTECH_XOR2 U140 ( .A(n164), .B(n139), .Z(n152) );
  GTECH_ADD_ABC U141 ( .A(n165), .B(n166), .C(n167), .COUT(n139) );
  GTECH_NOT U142 ( .A(n168), .Z(n167) );
  GTECH_XOR3 U143 ( .A(n169), .B(n170), .C(n171), .Z(n166) );
  GTECH_XOR4 U144 ( .A(n144), .B(n148), .C(n146), .D(n142), .Z(n164) );
  GTECH_XOR3 U145 ( .A(n134), .B(n136), .C(n135), .Z(n142) );
  GTECH_OAI21 U146 ( .A(n172), .B(n173), .C(n174), .Z(n135) );
  GTECH_OAI21 U147 ( .A(n175), .B(n176), .C(n177), .Z(n174) );
  GTECH_NOT U148 ( .A(n176), .Z(n172) );
  GTECH_NOT U149 ( .A(n178), .Z(n136) );
  GTECH_OR_NOT U150 ( .A(n179), .B(I_b[7]), .Z(n178) );
  GTECH_NOT U151 ( .A(n132), .Z(n134) );
  GTECH_OR_NOT U152 ( .A(n138), .B(I_b[6]), .Z(n132) );
  GTECH_NOT U153 ( .A(I_a[5]), .Z(n138) );
  GTECH_OR_NOT U154 ( .A(n180), .B(I_a[7]), .Z(n146) );
  GTECH_OAI21 U155 ( .A(n171), .B(n181), .C(n182), .Z(n148) );
  GTECH_OAI21 U156 ( .A(n169), .B(n183), .C(n170), .Z(n182) );
  GTECH_NOT U157 ( .A(n181), .Z(n169) );
  GTECH_NOT U158 ( .A(n183), .Z(n171) );
  GTECH_NOT U159 ( .A(n184), .Z(n144) );
  GTECH_OR_NOT U160 ( .A(n185), .B(I_a[6]), .Z(n184) );
  GTECH_OA22 U161 ( .A(n153), .B(n106), .C(n154), .D(n155), .Z(n159) );
  GTECH_NOT U162 ( .A(n186), .Z(n155) );
  GTECH_NOT U163 ( .A(I_a[7]), .Z(n106) );
  GTECH_XOR3 U164 ( .A(n156), .B(n161), .C(n187), .Z(N150) );
  GTECH_NOT U165 ( .A(n163), .Z(n187) );
  GTECH_XOR2 U166 ( .A(n188), .B(n165), .Z(n163) );
  GTECH_ADD_ABC U167 ( .A(n189), .B(n190), .C(n191), .COUT(n165) );
  GTECH_NOT U168 ( .A(n192), .Z(n191) );
  GTECH_XOR3 U169 ( .A(n193), .B(n194), .C(n195), .Z(n190) );
  GTECH_XOR4 U170 ( .A(n170), .B(n183), .C(n181), .D(n168), .Z(n188) );
  GTECH_XOR3 U171 ( .A(n175), .B(n177), .C(n176), .Z(n168) );
  GTECH_OAI21 U172 ( .A(n196), .B(n197), .C(n198), .Z(n176) );
  GTECH_OAI21 U173 ( .A(n199), .B(n200), .C(n201), .Z(n198) );
  GTECH_NOT U174 ( .A(n200), .Z(n196) );
  GTECH_NOT U175 ( .A(n202), .Z(n177) );
  GTECH_OR_NOT U176 ( .A(n203), .B(I_b[7]), .Z(n202) );
  GTECH_NOT U177 ( .A(n173), .Z(n175) );
  GTECH_OR_NOT U178 ( .A(n179), .B(I_b[6]), .Z(n173) );
  GTECH_OR_NOT U179 ( .A(n180), .B(I_a[6]), .Z(n181) );
  GTECH_OAI21 U180 ( .A(n195), .B(n204), .C(n205), .Z(n183) );
  GTECH_OAI21 U181 ( .A(n193), .B(n206), .C(n194), .Z(n205) );
  GTECH_NOT U182 ( .A(n204), .Z(n193) );
  GTECH_NOT U183 ( .A(n206), .Z(n195) );
  GTECH_NOT U184 ( .A(n207), .Z(n170) );
  GTECH_OR_NOT U185 ( .A(n185), .B(I_a[5]), .Z(n207) );
  GTECH_NOT U186 ( .A(I_b[5]), .Z(n185) );
  GTECH_NOT U187 ( .A(n157), .Z(n161) );
  GTECH_XOR2 U188 ( .A(n186), .B(n154), .Z(n157) );
  GTECH_AOI2N2 U189 ( .A(n208), .B(n209), .C(n210), .D(n211), .Z(n154) );
  GTECH_OR_NOT U190 ( .A(n212), .B(n210), .Z(n209) );
  GTECH_XOR2 U191 ( .A(n213), .B(n153), .Z(n186) );
  GTECH_AND2 U192 ( .A(n214), .B(n215), .Z(n153) );
  GTECH_OR_NOT U193 ( .A(n216), .B(n217), .Z(n215) );
  GTECH_OAI21 U194 ( .A(n218), .B(n217), .C(n219), .Z(n214) );
  GTECH_OR_NOT U195 ( .A(n220), .B(I_a[7]), .Z(n213) );
  GTECH_NOT U196 ( .A(n162), .Z(n156) );
  GTECH_OAI21 U197 ( .A(n221), .B(n222), .C(n223), .Z(n162) );
  GTECH_OAI21 U198 ( .A(n224), .B(n225), .C(n226), .Z(n223) );
  GTECH_NOT U199 ( .A(n221), .Z(n225) );
  GTECH_XOR3 U200 ( .A(n221), .B(n224), .C(n227), .Z(N149) );
  GTECH_NOT U201 ( .A(n226), .Z(n227) );
  GTECH_XOR2 U202 ( .A(n228), .B(n189), .Z(n226) );
  GTECH_ADD_ABC U203 ( .A(n229), .B(n230), .C(n231), .COUT(n189) );
  GTECH_XOR3 U204 ( .A(n232), .B(n233), .C(n234), .Z(n230) );
  GTECH_OA21 U205 ( .A(n235), .B(n236), .C(n237), .Z(n229) );
  GTECH_XOR4 U206 ( .A(n194), .B(n206), .C(n204), .D(n192), .Z(n228) );
  GTECH_XOR3 U207 ( .A(n199), .B(n201), .C(n200), .Z(n192) );
  GTECH_OAI21 U208 ( .A(n238), .B(n239), .C(n240), .Z(n200) );
  GTECH_NOT U209 ( .A(n241), .Z(n201) );
  GTECH_OR_NOT U210 ( .A(n242), .B(I_b[7]), .Z(n241) );
  GTECH_NOT U211 ( .A(n197), .Z(n199) );
  GTECH_OR_NOT U212 ( .A(n203), .B(I_b[6]), .Z(n197) );
  GTECH_OR_NOT U213 ( .A(n180), .B(I_a[5]), .Z(n204) );
  GTECH_NOT U214 ( .A(I_b[4]), .Z(n180) );
  GTECH_OAI21 U215 ( .A(n234), .B(n243), .C(n244), .Z(n206) );
  GTECH_OAI21 U216 ( .A(n232), .B(n245), .C(n233), .Z(n244) );
  GTECH_NOT U217 ( .A(n243), .Z(n232) );
  GTECH_NOT U218 ( .A(n245), .Z(n234) );
  GTECH_NOT U219 ( .A(n246), .Z(n194) );
  GTECH_OR_NOT U220 ( .A(n179), .B(I_b[5]), .Z(n246) );
  GTECH_NOT U221 ( .A(n222), .Z(n224) );
  GTECH_XOR3 U222 ( .A(n212), .B(n210), .C(n208), .Z(n222) );
  GTECH_XOR3 U223 ( .A(n218), .B(n219), .C(n217), .Z(n208) );
  GTECH_OAI21 U224 ( .A(n247), .B(n248), .C(n249), .Z(n217) );
  GTECH_OAI21 U225 ( .A(n250), .B(n251), .C(n252), .Z(n249) );
  GTECH_NOT U226 ( .A(n251), .Z(n247) );
  GTECH_NOT U227 ( .A(n253), .Z(n219) );
  GTECH_OR_NOT U228 ( .A(n220), .B(I_a[6]), .Z(n253) );
  GTECH_NOT U229 ( .A(n216), .Z(n218) );
  GTECH_OR_NOT U230 ( .A(n254), .B(I_a[7]), .Z(n216) );
  GTECH_ADD_ABC U231 ( .A(n255), .B(n256), .C(n257), .COUT(n210) );
  GTECH_XOR2 U232 ( .A(n258), .B(n259), .Z(n256) );
  GTECH_AND2 U233 ( .A(I_a[7]), .B(I_b[1]), .Z(n259) );
  GTECH_NOT U234 ( .A(n211), .Z(n212) );
  GTECH_OR_NOT U235 ( .A(n258), .B(I_a[7]), .Z(n211) );
  GTECH_ADD_ABC U236 ( .A(n260), .B(n261), .C(n262), .COUT(n221) );
  GTECH_XOR3 U237 ( .A(n255), .B(n263), .C(n257), .Z(n261) );
  GTECH_NOT U238 ( .A(n264), .Z(n257) );
  GTECH_XOR2 U239 ( .A(n260), .B(n265), .Z(N148) );
  GTECH_XOR4 U240 ( .A(n263), .B(n264), .C(n262), .D(n255), .Z(n265) );
  GTECH_ADD_ABC U241 ( .A(n266), .B(n267), .C(n268), .COUT(n255) );
  GTECH_XOR3 U242 ( .A(n269), .B(n270), .C(n271), .Z(n267) );
  GTECH_XOR2 U243 ( .A(n272), .B(n273), .Z(n262) );
  GTECH_OA21 U244 ( .A(n235), .B(n236), .C(n237), .Z(n273) );
  GTECH_OAI21 U245 ( .A(n274), .B(n275), .C(n276), .Z(n237) );
  GTECH_NOT U246 ( .A(n235), .Z(n275) );
  GTECH_XOR4 U247 ( .A(n233), .B(n245), .C(n243), .D(n231), .Z(n272) );
  GTECH_XOR3 U248 ( .A(n277), .B(n278), .C(n240), .Z(n231) );
  GTECH_NAND3 U249 ( .A(I_b[6]), .B(I_a[1]), .C(n279), .Z(n240) );
  GTECH_NOT U250 ( .A(n239), .Z(n278) );
  GTECH_OR_NOT U251 ( .A(n280), .B(I_b[7]), .Z(n239) );
  GTECH_NOT U252 ( .A(n238), .Z(n277) );
  GTECH_OR_NOT U253 ( .A(n242), .B(I_b[6]), .Z(n238) );
  GTECH_OR_NOT U254 ( .A(n179), .B(I_b[4]), .Z(n243) );
  GTECH_OAI21 U255 ( .A(n281), .B(n282), .C(n283), .Z(n245) );
  GTECH_OAI21 U256 ( .A(n284), .B(n285), .C(n286), .Z(n283) );
  GTECH_NOT U257 ( .A(n285), .Z(n281) );
  GTECH_NOT U258 ( .A(n287), .Z(n233) );
  GTECH_OR_NOT U259 ( .A(n203), .B(I_b[5]), .Z(n287) );
  GTECH_XOR3 U260 ( .A(n250), .B(n252), .C(n251), .Z(n264) );
  GTECH_OAI21 U261 ( .A(n288), .B(n289), .C(n290), .Z(n251) );
  GTECH_OAI21 U262 ( .A(n291), .B(n292), .C(n293), .Z(n290) );
  GTECH_NOT U263 ( .A(n292), .Z(n288) );
  GTECH_NOT U264 ( .A(n294), .Z(n252) );
  GTECH_OR_NOT U265 ( .A(n220), .B(I_a[5]), .Z(n294) );
  GTECH_NOT U266 ( .A(I_b[3]), .Z(n220) );
  GTECH_NOT U267 ( .A(n248), .Z(n250) );
  GTECH_OR_NOT U268 ( .A(n254), .B(I_a[6]), .Z(n248) );
  GTECH_XOR2 U269 ( .A(n295), .B(n258), .Z(n263) );
  GTECH_OA21 U270 ( .A(n271), .B(n296), .C(n297), .Z(n258) );
  GTECH_OAI21 U271 ( .A(n269), .B(n298), .C(n270), .Z(n297) );
  GTECH_NOT U272 ( .A(n298), .Z(n271) );
  GTECH_AND2 U273 ( .A(I_b[1]), .B(I_a[7]), .Z(n295) );
  GTECH_ADD_ABC U274 ( .A(n299), .B(n300), .C(n301), .COUT(n260) );
  GTECH_NOT U275 ( .A(n302), .Z(n301) );
  GTECH_XOR3 U276 ( .A(n266), .B(n303), .C(n268), .Z(n300) );
  GTECH_NOT U277 ( .A(n304), .Z(n268) );
  GTECH_NOT U278 ( .A(n305), .Z(n303) );
  GTECH_XOR2 U279 ( .A(n306), .B(n299), .Z(N147) );
  GTECH_ADD_ABC U280 ( .A(n307), .B(n308), .C(n309), .COUT(n299) );
  GTECH_XOR3 U281 ( .A(n310), .B(n311), .C(n312), .Z(n308) );
  GTECH_OA21 U282 ( .A(n313), .B(n314), .C(n315), .Z(n307) );
  GTECH_XOR4 U283 ( .A(n304), .B(n266), .C(n305), .D(n302), .Z(n306) );
  GTECH_XOR3 U284 ( .A(n276), .B(n236), .C(n235), .Z(n302) );
  GTECH_XOR2 U285 ( .A(n316), .B(n279), .Z(n235) );
  GTECH_NOT U286 ( .A(n317), .Z(n279) );
  GTECH_OR_NOT U287 ( .A(n318), .B(I_b[7]), .Z(n317) );
  GTECH_OR_NOT U288 ( .A(n280), .B(I_b[6]), .Z(n316) );
  GTECH_NOT U289 ( .A(n274), .Z(n236) );
  GTECH_XOR3 U290 ( .A(n284), .B(n286), .C(n285), .Z(n274) );
  GTECH_OAI21 U291 ( .A(n319), .B(n320), .C(n321), .Z(n285) );
  GTECH_NOT U292 ( .A(n322), .Z(n286) );
  GTECH_OR_NOT U293 ( .A(n242), .B(I_b[5]), .Z(n322) );
  GTECH_NOT U294 ( .A(n282), .Z(n284) );
  GTECH_OR_NOT U295 ( .A(n203), .B(I_b[4]), .Z(n282) );
  GTECH_NOT U296 ( .A(n323), .Z(n276) );
  GTECH_NAND3 U297 ( .A(I_a[0]), .B(n324), .C(I_b[6]), .Z(n323) );
  GTECH_NOT U298 ( .A(n325), .Z(n324) );
  GTECH_XOR3 U299 ( .A(n269), .B(n270), .C(n298), .Z(n305) );
  GTECH_OAI21 U300 ( .A(n326), .B(n327), .C(n328), .Z(n298) );
  GTECH_OAI21 U301 ( .A(n329), .B(n330), .C(n331), .Z(n328) );
  GTECH_NOT U302 ( .A(n332), .Z(n270) );
  GTECH_OR_NOT U303 ( .A(n333), .B(I_a[6]), .Z(n332) );
  GTECH_NOT U304 ( .A(n296), .Z(n269) );
  GTECH_OR_NOT U305 ( .A(n334), .B(I_a[7]), .Z(n296) );
  GTECH_ADD_ABC U306 ( .A(n310), .B(n335), .C(n312), .COUT(n266) );
  GTECH_NOT U307 ( .A(n336), .Z(n312) );
  GTECH_XOR3 U308 ( .A(n329), .B(n331), .C(n326), .Z(n335) );
  GTECH_NOT U309 ( .A(n330), .Z(n326) );
  GTECH_XOR3 U310 ( .A(n291), .B(n293), .C(n292), .Z(n304) );
  GTECH_OAI21 U311 ( .A(n337), .B(n338), .C(n339), .Z(n292) );
  GTECH_OAI21 U312 ( .A(n340), .B(n341), .C(n342), .Z(n339) );
  GTECH_NOT U313 ( .A(n341), .Z(n337) );
  GTECH_NOT U314 ( .A(n343), .Z(n293) );
  GTECH_OR_NOT U315 ( .A(n179), .B(I_b[3]), .Z(n343) );
  GTECH_NOT U316 ( .A(n289), .Z(n291) );
  GTECH_OR_NOT U317 ( .A(n254), .B(I_a[5]), .Z(n289) );
  GTECH_NOT U318 ( .A(I_b[2]), .Z(n254) );
  GTECH_XOR2 U319 ( .A(n344), .B(n345), .Z(N146) );
  GTECH_XOR4 U320 ( .A(n311), .B(n336), .C(n309), .D(n310), .Z(n345) );
  GTECH_ADD_ABC U321 ( .A(n346), .B(n347), .C(n348), .COUT(n310) );
  GTECH_NOT U322 ( .A(n349), .Z(n348) );
  GTECH_XOR3 U323 ( .A(n350), .B(n351), .C(n352), .Z(n347) );
  GTECH_XOR2 U324 ( .A(n325), .B(n353), .Z(n309) );
  GTECH_AND2 U325 ( .A(I_b[6]), .B(I_a[0]), .Z(n353) );
  GTECH_XOR3 U326 ( .A(n354), .B(n355), .C(n321), .Z(n325) );
  GTECH_NAND3 U327 ( .A(I_b[4]), .B(I_a[1]), .C(n356), .Z(n321) );
  GTECH_NOT U328 ( .A(n320), .Z(n355) );
  GTECH_OR_NOT U329 ( .A(n280), .B(I_b[5]), .Z(n320) );
  GTECH_NOT U330 ( .A(n319), .Z(n354) );
  GTECH_OR_NOT U331 ( .A(n242), .B(I_b[4]), .Z(n319) );
  GTECH_XOR3 U332 ( .A(n340), .B(n342), .C(n341), .Z(n336) );
  GTECH_OAI21 U333 ( .A(n357), .B(n358), .C(n359), .Z(n341) );
  GTECH_OAI21 U334 ( .A(n360), .B(n361), .C(n362), .Z(n359) );
  GTECH_NOT U335 ( .A(n361), .Z(n357) );
  GTECH_NOT U336 ( .A(n363), .Z(n342) );
  GTECH_OR_NOT U337 ( .A(n203), .B(I_b[3]), .Z(n363) );
  GTECH_NOT U338 ( .A(n338), .Z(n340) );
  GTECH_OR_NOT U339 ( .A(n179), .B(I_b[2]), .Z(n338) );
  GTECH_NOT U340 ( .A(I_a[4]), .Z(n179) );
  GTECH_NOT U341 ( .A(n364), .Z(n311) );
  GTECH_XOR3 U342 ( .A(n329), .B(n331), .C(n330), .Z(n364) );
  GTECH_OAI21 U343 ( .A(n352), .B(n365), .C(n366), .Z(n330) );
  GTECH_OAI21 U344 ( .A(n350), .B(n367), .C(n351), .Z(n366) );
  GTECH_NOT U345 ( .A(n365), .Z(n350) );
  GTECH_NOT U346 ( .A(n367), .Z(n352) );
  GTECH_NOT U347 ( .A(n368), .Z(n331) );
  GTECH_OR_NOT U348 ( .A(n333), .B(I_a[5]), .Z(n368) );
  GTECH_NOT U349 ( .A(n327), .Z(n329) );
  GTECH_OR_NOT U350 ( .A(n334), .B(I_a[6]), .Z(n327) );
  GTECH_OA21 U351 ( .A(n313), .B(n314), .C(n315), .Z(n344) );
  GTECH_OAI21 U352 ( .A(n369), .B(n370), .C(n371), .Z(n315) );
  GTECH_NOT U353 ( .A(n313), .Z(n370) );
  GTECH_XOR3 U354 ( .A(n371), .B(n314), .C(n313), .Z(N145) );
  GTECH_XOR2 U355 ( .A(n372), .B(n356), .Z(n313) );
  GTECH_NOT U356 ( .A(n373), .Z(n356) );
  GTECH_OR_NOT U357 ( .A(n318), .B(I_b[5]), .Z(n373) );
  GTECH_OR_NOT U358 ( .A(n280), .B(I_b[4]), .Z(n372) );
  GTECH_NOT U359 ( .A(n369), .Z(n314) );
  GTECH_XOR2 U360 ( .A(n374), .B(n346), .Z(n369) );
  GTECH_ADD_ABC U361 ( .A(n375), .B(n376), .C(n377), .COUT(n346) );
  GTECH_XOR3 U362 ( .A(n378), .B(n379), .C(n380), .Z(n376) );
  GTECH_OA21 U363 ( .A(n381), .B(n382), .C(n383), .Z(n375) );
  GTECH_XOR4 U364 ( .A(n351), .B(n367), .C(n365), .D(n349), .Z(n374) );
  GTECH_XOR3 U365 ( .A(n360), .B(n362), .C(n361), .Z(n349) );
  GTECH_OAI21 U366 ( .A(n384), .B(n385), .C(n386), .Z(n361) );
  GTECH_NOT U367 ( .A(n387), .Z(n362) );
  GTECH_OR_NOT U368 ( .A(n242), .B(I_b[3]), .Z(n387) );
  GTECH_NOT U369 ( .A(n358), .Z(n360) );
  GTECH_OR_NOT U370 ( .A(n203), .B(I_b[2]), .Z(n358) );
  GTECH_OR_NOT U371 ( .A(n334), .B(I_a[5]), .Z(n365) );
  GTECH_OAI21 U372 ( .A(n380), .B(n388), .C(n389), .Z(n367) );
  GTECH_OAI21 U373 ( .A(n378), .B(n390), .C(n379), .Z(n389) );
  GTECH_NOT U374 ( .A(n390), .Z(n380) );
  GTECH_NOT U375 ( .A(n391), .Z(n351) );
  GTECH_OR_NOT U376 ( .A(n333), .B(I_a[4]), .Z(n391) );
  GTECH_NOT U377 ( .A(n392), .Z(n371) );
  GTECH_NAND3 U378 ( .A(I_a[0]), .B(n393), .C(I_b[4]), .Z(n392) );
  GTECH_XOR2 U379 ( .A(n394), .B(n393), .Z(N144) );
  GTECH_XOR2 U380 ( .A(n395), .B(n396), .Z(n393) );
  GTECH_XOR4 U381 ( .A(n379), .B(n390), .C(n377), .D(n378), .Z(n396) );
  GTECH_NOT U382 ( .A(n388), .Z(n378) );
  GTECH_OR_NOT U383 ( .A(n334), .B(I_a[4]), .Z(n388) );
  GTECH_NOT U384 ( .A(I_b[0]), .Z(n334) );
  GTECH_XOR3 U385 ( .A(n397), .B(n398), .C(n386), .Z(n377) );
  GTECH_NAND3 U386 ( .A(I_b[2]), .B(I_a[1]), .C(n399), .Z(n386) );
  GTECH_NOT U387 ( .A(n385), .Z(n398) );
  GTECH_OR_NOT U388 ( .A(n280), .B(I_b[3]), .Z(n385) );
  GTECH_NOT U389 ( .A(n384), .Z(n397) );
  GTECH_OR_NOT U390 ( .A(n242), .B(I_b[2]), .Z(n384) );
  GTECH_OAI21 U391 ( .A(n400), .B(n401), .C(n402), .Z(n390) );
  GTECH_OAI21 U392 ( .A(n403), .B(n404), .C(n405), .Z(n402) );
  GTECH_NOT U393 ( .A(n404), .Z(n400) );
  GTECH_NOT U394 ( .A(n406), .Z(n379) );
  GTECH_OR_NOT U395 ( .A(n333), .B(I_a[3]), .Z(n406) );
  GTECH_OA21 U396 ( .A(n381), .B(n382), .C(n383), .Z(n395) );
  GTECH_OAI21 U397 ( .A(n407), .B(n408), .C(n409), .Z(n383) );
  GTECH_NOT U398 ( .A(n381), .Z(n408) );
  GTECH_AND2 U399 ( .A(I_b[4]), .B(I_a[0]), .Z(n394) );
  GTECH_XOR3 U400 ( .A(n409), .B(n382), .C(n381), .Z(N143) );
  GTECH_XOR2 U401 ( .A(n410), .B(n399), .Z(n381) );
  GTECH_NOT U402 ( .A(n411), .Z(n399) );
  GTECH_OR_NOT U403 ( .A(n318), .B(I_b[3]), .Z(n411) );
  GTECH_NOT U404 ( .A(I_a[0]), .Z(n318) );
  GTECH_OR_NOT U405 ( .A(n280), .B(I_b[2]), .Z(n410) );
  GTECH_NOT U406 ( .A(I_a[1]), .Z(n280) );
  GTECH_NOT U407 ( .A(n407), .Z(n382) );
  GTECH_XOR3 U408 ( .A(n403), .B(n405), .C(n404), .Z(n407) );
  GTECH_OAI21 U409 ( .A(n412), .B(n413), .C(n414), .Z(n404) );
  GTECH_NOT U410 ( .A(n415), .Z(n405) );
  GTECH_OR_NOT U411 ( .A(n242), .B(I_b[1]), .Z(n415) );
  GTECH_NOT U412 ( .A(n401), .Z(n403) );
  GTECH_OR_NOT U413 ( .A(n203), .B(I_b[0]), .Z(n401) );
  GTECH_NOT U414 ( .A(I_a[3]), .Z(n203) );
  GTECH_NOT U415 ( .A(n416), .Z(n409) );
  GTECH_NAND3 U416 ( .A(I_a[0]), .B(n417), .C(I_b[2]), .Z(n416) );
  GTECH_XOR2 U417 ( .A(n418), .B(n417), .Z(N142) );
  GTECH_NOT U418 ( .A(n419), .Z(n417) );
  GTECH_XOR3 U419 ( .A(n420), .B(n421), .C(n414), .Z(n419) );
  GTECH_NAND3 U420 ( .A(n422), .B(I_b[0]), .C(I_a[1]), .Z(n414) );
  GTECH_NOT U421 ( .A(n412), .Z(n421) );
  GTECH_OR_NOT U422 ( .A(n333), .B(I_a[1]), .Z(n412) );
  GTECH_NOT U423 ( .A(n413), .Z(n420) );
  GTECH_OR_NOT U424 ( .A(n242), .B(I_b[0]), .Z(n413) );
  GTECH_NOT U425 ( .A(I_a[2]), .Z(n242) );
  GTECH_AND2 U426 ( .A(I_b[2]), .B(I_a[0]), .Z(n418) );
  GTECH_XOR2 U427 ( .A(n422), .B(n423), .Z(N141) );
  GTECH_AND2 U428 ( .A(I_a[1]), .B(I_b[0]), .Z(n423) );
  GTECH_NOT U429 ( .A(n424), .Z(n422) );
  GTECH_OR_NOT U430 ( .A(n333), .B(I_a[0]), .Z(n424) );
  GTECH_NOT U431 ( .A(I_b[1]), .Z(n333) );
  GTECH_AND2 U432 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

