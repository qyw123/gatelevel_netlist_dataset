
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385;

  GTECH_MUX2 U137 ( .A(n276), .B(n277), .S(n278), .Z(sum[9]) );
  GTECH_XOR2 U138 ( .A(n279), .B(n280), .Z(n277) );
  GTECH_XOR2 U139 ( .A(n281), .B(n280), .Z(n276) );
  GTECH_OA21 U140 ( .A(b[9]), .B(a[9]), .C(n282), .Z(n280) );
  GTECH_NOT U141 ( .A(n283), .Z(n282) );
  GTECH_XNOR2 U142 ( .A(n278), .B(n284), .Z(sum[8]) );
  GTECH_MUX2 U143 ( .A(n285), .B(n286), .S(n287), .Z(sum[7]) );
  GTECH_XOR2 U144 ( .A(n288), .B(n289), .Z(n286) );
  GTECH_XNOR2 U145 ( .A(n288), .B(n290), .Z(n285) );
  GTECH_NOR2 U146 ( .A(n291), .B(n292), .Z(n290) );
  GTECH_OA21 U147 ( .A(a[6]), .B(b[6]), .C(n293), .Z(n292) );
  GTECH_XOR2 U148 ( .A(a[7]), .B(b[7]), .Z(n288) );
  GTECH_AO21 U149 ( .A(n291), .B(n294), .C(n295), .Z(sum[6]) );
  GTECH_MUX2 U150 ( .A(n296), .B(n297), .S(b[6]), .Z(n295) );
  GTECH_AND2 U151 ( .A(n298), .B(n299), .Z(n297) );
  GTECH_XNOR2 U152 ( .A(a[6]), .B(n298), .Z(n296) );
  GTECH_NOT U153 ( .A(n294), .Z(n298) );
  GTECH_OA21 U154 ( .A(n287), .B(n293), .C(n300), .Z(n294) );
  GTECH_OA21 U155 ( .A(n301), .B(n302), .C(n303), .Z(n293) );
  GTECH_MUX2 U156 ( .A(n304), .B(n305), .S(n306), .Z(sum[5]) );
  GTECH_AND_NOT U157 ( .A(n303), .B(n301), .Z(n306) );
  GTECH_NOT U158 ( .A(n307), .Z(n305) );
  GTECH_OA21 U159 ( .A(n287), .B(n302), .C(n308), .Z(n307) );
  GTECH_AO21 U160 ( .A(n287), .B(n308), .C(n302), .Z(n304) );
  GTECH_XOR2 U161 ( .A(n309), .B(n287), .Z(sum[4]) );
  GTECH_MUX2 U162 ( .A(n310), .B(n311), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U163 ( .A(n312), .B(n313), .Z(n311) );
  GTECH_XNOR2 U164 ( .A(n312), .B(n314), .Z(n310) );
  GTECH_NOR2 U165 ( .A(n315), .B(n316), .Z(n314) );
  GTECH_OA21 U166 ( .A(a[2]), .B(b[2]), .C(n317), .Z(n316) );
  GTECH_XOR2 U167 ( .A(a[3]), .B(b[3]), .Z(n312) );
  GTECH_MUX2 U168 ( .A(n318), .B(n319), .S(cin), .Z(sum[2]) );
  GTECH_MUX2 U169 ( .A(n320), .B(n321), .S(n322), .Z(n319) );
  GTECH_MUX2 U170 ( .A(n320), .B(n321), .S(n317), .Z(n318) );
  GTECH_OA21 U171 ( .A(n323), .B(n324), .C(n325), .Z(n317) );
  GTECH_AO21 U172 ( .A(n326), .B(n327), .C(n315), .Z(n321) );
  GTECH_XNOR2 U173 ( .A(a[2]), .B(n327), .Z(n320) );
  GTECH_NOT U174 ( .A(b[2]), .Z(n327) );
  GTECH_MUX2 U175 ( .A(n328), .B(n329), .S(n330), .Z(sum[1]) );
  GTECH_AND_NOT U176 ( .A(n325), .B(n324), .Z(n330) );
  GTECH_NOT U177 ( .A(n331), .Z(n329) );
  GTECH_OA21 U178 ( .A(n323), .B(cin), .C(n332), .Z(n331) );
  GTECH_AO21 U179 ( .A(cin), .B(n332), .C(n323), .Z(n328) );
  GTECH_AND2 U180 ( .A(a[0]), .B(b[0]), .Z(n323) );
  GTECH_MUX2 U181 ( .A(n333), .B(n334), .S(n335), .Z(sum[15]) );
  GTECH_XNOR2 U182 ( .A(n336), .B(n337), .Z(n334) );
  GTECH_AND_NOT U183 ( .A(n338), .B(n339), .Z(n337) );
  GTECH_AO21 U184 ( .A(n340), .B(n341), .C(n342), .Z(n338) );
  GTECH_XOR2 U185 ( .A(n336), .B(n343), .Z(n333) );
  GTECH_XOR2 U186 ( .A(a[15]), .B(b[15]), .Z(n336) );
  GTECH_AO21 U187 ( .A(n339), .B(n344), .C(n345), .Z(sum[14]) );
  GTECH_MUX2 U188 ( .A(n346), .B(n347), .S(n341), .Z(n345) );
  GTECH_XNOR2 U189 ( .A(a[14]), .B(n348), .Z(n347) );
  GTECH_AND2 U190 ( .A(n348), .B(n340), .Z(n346) );
  GTECH_NOT U191 ( .A(n348), .Z(n344) );
  GTECH_AO21 U192 ( .A(n335), .B(n342), .C(n349), .Z(n348) );
  GTECH_OAI22 U193 ( .A(b[13]), .B(a[13]), .C(n350), .D(n351), .Z(n342) );
  GTECH_MUX2 U194 ( .A(n352), .B(n353), .S(n335), .Z(sum[13]) );
  GTECH_MUX2 U195 ( .A(n354), .B(n355), .S(n351), .Z(n353) );
  GTECH_MUX2 U196 ( .A(n354), .B(n355), .S(n356), .Z(n352) );
  GTECH_AO21 U197 ( .A(n357), .B(n358), .C(n350), .Z(n355) );
  GTECH_XNOR2 U198 ( .A(a[13]), .B(n357), .Z(n354) );
  GTECH_NOT U199 ( .A(b[13]), .Z(n357) );
  GTECH_XNOR2 U200 ( .A(n359), .B(n335), .Z(sum[12]) );
  GTECH_MUX2 U201 ( .A(n360), .B(n361), .S(n278), .Z(sum[11]) );
  GTECH_XOR2 U202 ( .A(n362), .B(n363), .Z(n361) );
  GTECH_XNOR2 U203 ( .A(n362), .B(n364), .Z(n360) );
  GTECH_AOI21 U204 ( .A(n365), .B(n366), .C(n367), .Z(n364) );
  GTECH_XOR2 U205 ( .A(a[11]), .B(b[11]), .Z(n362) );
  GTECH_MUX2 U206 ( .A(n368), .B(n369), .S(n278), .Z(sum[10]) );
  GTECH_XNOR2 U207 ( .A(n370), .B(n371), .Z(n369) );
  GTECH_XNOR2 U208 ( .A(n370), .B(n366), .Z(n368) );
  GTECH_OA21 U209 ( .A(n283), .B(n281), .C(n372), .Z(n366) );
  GTECH_OR_NOT U210 ( .A(n367), .B(n365), .Z(n370) );
  GTECH_XNOR2 U211 ( .A(cin), .B(n373), .Z(sum[0]) );
  GTECH_MUX2 U212 ( .A(n374), .B(n359), .S(n335), .Z(cout) );
  GTECH_MUX2 U213 ( .A(n284), .B(n375), .S(n278), .Z(n335) );
  GTECH_MUX2 U214 ( .A(n309), .B(n376), .S(n287), .Z(n278) );
  GTECH_NOT U215 ( .A(n377), .Z(n287) );
  GTECH_MUX2 U216 ( .A(n373), .B(n378), .S(cin), .Z(n377) );
  GTECH_AOI21 U217 ( .A(n313), .B(a[3]), .C(n379), .Z(n378) );
  GTECH_OA21 U218 ( .A(n313), .B(a[3]), .C(b[3]), .Z(n379) );
  GTECH_OR2 U219 ( .A(n380), .B(n315), .Z(n313) );
  GTECH_AND_NOT U220 ( .A(b[2]), .B(n326), .Z(n315) );
  GTECH_NOT U221 ( .A(a[2]), .Z(n326) );
  GTECH_OA21 U222 ( .A(b[2]), .B(a[2]), .C(n322), .Z(n380) );
  GTECH_OA21 U223 ( .A(n332), .B(n324), .C(n325), .Z(n322) );
  GTECH_OR2 U224 ( .A(a[1]), .B(b[1]), .Z(n325) );
  GTECH_AND2 U225 ( .A(a[1]), .B(b[1]), .Z(n324) );
  GTECH_OR2 U226 ( .A(a[0]), .B(b[0]), .Z(n332) );
  GTECH_XNOR2 U227 ( .A(a[0]), .B(b[0]), .Z(n373) );
  GTECH_OA21 U228 ( .A(a[7]), .B(n289), .C(n381), .Z(n376) );
  GTECH_AO21 U229 ( .A(a[7]), .B(n289), .C(b[7]), .Z(n381) );
  GTECH_OR2 U230 ( .A(n382), .B(n291), .Z(n289) );
  GTECH_AND_NOT U231 ( .A(b[6]), .B(n299), .Z(n291) );
  GTECH_NOT U232 ( .A(a[6]), .Z(n299) );
  GTECH_OA21 U233 ( .A(b[6]), .B(a[6]), .C(n300), .Z(n382) );
  GTECH_OA21 U234 ( .A(n308), .B(n301), .C(n303), .Z(n300) );
  GTECH_OR2 U235 ( .A(a[5]), .B(b[5]), .Z(n303) );
  GTECH_AND2 U236 ( .A(a[5]), .B(b[5]), .Z(n301) );
  GTECH_AND_NOT U237 ( .A(n308), .B(n302), .Z(n309) );
  GTECH_AND2 U238 ( .A(b[4]), .B(a[4]), .Z(n302) );
  GTECH_OR2 U239 ( .A(b[4]), .B(a[4]), .Z(n308) );
  GTECH_AOI21 U240 ( .A(n363), .B(a[11]), .C(n383), .Z(n375) );
  GTECH_OA21 U241 ( .A(n363), .B(a[11]), .C(b[11]), .Z(n383) );
  GTECH_AO21 U242 ( .A(n371), .B(n365), .C(n367), .Z(n363) );
  GTECH_AND2 U243 ( .A(b[10]), .B(a[10]), .Z(n367) );
  GTECH_OR2 U244 ( .A(a[10]), .B(b[10]), .Z(n365) );
  GTECH_OA21 U245 ( .A(n279), .B(n283), .C(n372), .Z(n371) );
  GTECH_OR2 U246 ( .A(a[9]), .B(b[9]), .Z(n372) );
  GTECH_AND2 U247 ( .A(a[9]), .B(b[9]), .Z(n283) );
  GTECH_OR_NOT U248 ( .A(n281), .B(n279), .Z(n284) );
  GTECH_OR2 U249 ( .A(b[8]), .B(a[8]), .Z(n279) );
  GTECH_AND2 U250 ( .A(a[8]), .B(b[8]), .Z(n281) );
  GTECH_AND_NOT U251 ( .A(n356), .B(n351), .Z(n359) );
  GTECH_AND2 U252 ( .A(a[12]), .B(b[12]), .Z(n351) );
  GTECH_AO22 U253 ( .A(n384), .B(b[15]), .C(n343), .D(a[15]), .Z(n374) );
  GTECH_OR2 U254 ( .A(n343), .B(a[15]), .Z(n384) );
  GTECH_OR_NOT U255 ( .A(n339), .B(n385), .Z(n343) );
  GTECH_AO21 U256 ( .A(n341), .B(n340), .C(n349), .Z(n385) );
  GTECH_OAI22 U257 ( .A(n350), .B(n356), .C(b[13]), .D(a[13]), .Z(n349) );
  GTECH_OR2 U258 ( .A(a[12]), .B(b[12]), .Z(n356) );
  GTECH_AND_NOT U259 ( .A(b[13]), .B(n358), .Z(n350) );
  GTECH_NOT U260 ( .A(a[13]), .Z(n358) );
  GTECH_NOT U261 ( .A(b[14]), .Z(n341) );
  GTECH_AND_NOT U262 ( .A(b[14]), .B(n340), .Z(n339) );
  GTECH_NOT U263 ( .A(a[14]), .Z(n340) );
endmodule

