
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394;

  GTECH_MUX2 U137 ( .A(n276), .B(n277), .S(n278), .Z(sum[9]) );
  GTECH_OA21 U138 ( .A(n279), .B(n280), .C(n281), .Z(n278) );
  GTECH_OAI21 U139 ( .A(a[8]), .B(n282), .C(b[8]), .Z(n281) );
  GTECH_NOT U140 ( .A(n282), .Z(n279) );
  GTECH_XOR2 U141 ( .A(b[9]), .B(a[9]), .Z(n277) );
  GTECH_OR2 U142 ( .A(n283), .B(n284), .Z(n276) );
  GTECH_AO21 U143 ( .A(n282), .B(n285), .C(n286), .Z(sum[8]) );
  GTECH_MUX2 U144 ( .A(n287), .B(n288), .S(n289), .Z(sum[7]) );
  GTECH_XOR2 U145 ( .A(n290), .B(n291), .Z(n288) );
  GTECH_XOR2 U146 ( .A(n292), .B(n290), .Z(n287) );
  GTECH_XOR2 U147 ( .A(a[7]), .B(b[7]), .Z(n290) );
  GTECH_OA21 U148 ( .A(a[6]), .B(n293), .C(n294), .Z(n292) );
  GTECH_AO21 U149 ( .A(n293), .B(a[6]), .C(b[6]), .Z(n294) );
  GTECH_MUX2 U150 ( .A(n295), .B(n296), .S(n289), .Z(sum[6]) );
  GTECH_XOR2 U151 ( .A(n297), .B(n298), .Z(n296) );
  GTECH_XOR2 U152 ( .A(n297), .B(n293), .Z(n295) );
  GTECH_AO21 U153 ( .A(a[4]), .B(n299), .C(n300), .Z(n293) );
  GTECH_AND_NOT U154 ( .A(b[4]), .B(n301), .Z(n299) );
  GTECH_XOR2 U155 ( .A(a[6]), .B(b[6]), .Z(n297) );
  GTECH_XOR2 U156 ( .A(n302), .B(n303), .Z(sum[5]) );
  GTECH_ADD_ABC U157 ( .A(a[4]), .B(n304), .C(b[4]), .COUT(n303) );
  GTECH_MUX2 U158 ( .A(n305), .B(n306), .S(n307), .Z(n304) );
  GTECH_OAI21 U159 ( .A(n308), .B(n309), .C(n310), .Z(n305) );
  GTECH_NOR2 U160 ( .A(n300), .B(n301), .Z(n302) );
  GTECH_XOR2 U161 ( .A(n289), .B(n311), .Z(sum[4]) );
  GTECH_MUX2 U162 ( .A(n312), .B(n313), .S(n307), .Z(sum[3]) );
  GTECH_XOR2 U163 ( .A(n314), .B(n315), .Z(n313) );
  GTECH_OAI21 U164 ( .A(a[2]), .B(n316), .C(n317), .Z(n314) );
  GTECH_AO21 U165 ( .A(n316), .B(a[2]), .C(b[2]), .Z(n317) );
  GTECH_XOR2 U166 ( .A(n315), .B(n308), .Z(n312) );
  GTECH_XOR2 U167 ( .A(n309), .B(b[3]), .Z(n315) );
  GTECH_MUX2 U168 ( .A(n318), .B(n319), .S(n307), .Z(sum[2]) );
  GTECH_XOR2 U169 ( .A(n320), .B(n316), .Z(n319) );
  GTECH_ADD_ABC U170 ( .A(a[1]), .B(n321), .C(b[1]), .COUT(n316) );
  GTECH_AND2 U171 ( .A(a[0]), .B(b[0]), .Z(n321) );
  GTECH_XOR2 U172 ( .A(n322), .B(n320), .Z(n318) );
  GTECH_XOR2 U173 ( .A(a[2]), .B(b[2]), .Z(n320) );
  GTECH_MUX2 U174 ( .A(n323), .B(n324), .S(n325), .Z(sum[1]) );
  GTECH_XOR2 U175 ( .A(b[1]), .B(a[1]), .Z(n325) );
  GTECH_AO21 U176 ( .A(n307), .B(n326), .C(n327), .Z(n324) );
  GTECH_OAI21 U177 ( .A(n327), .B(n307), .C(n326), .Z(n323) );
  GTECH_OR_NOT U178 ( .A(n328), .B(a[0]), .Z(n326) );
  GTECH_MUX2 U179 ( .A(n329), .B(n330), .S(n331), .Z(sum[15]) );
  GTECH_XOR2 U180 ( .A(n332), .B(n333), .Z(n330) );
  GTECH_XOR2 U181 ( .A(n332), .B(n334), .Z(n329) );
  GTECH_AND_NOT U182 ( .A(n335), .B(n336), .Z(n334) );
  GTECH_OAI21 U183 ( .A(b[14]), .B(a[14]), .C(n337), .Z(n335) );
  GTECH_XOR2 U184 ( .A(n338), .B(b[15]), .Z(n332) );
  GTECH_MUX2 U185 ( .A(n339), .B(n340), .S(n341), .Z(sum[14]) );
  GTECH_XOR2 U186 ( .A(n342), .B(n337), .Z(n340) );
  GTECH_OAI21 U187 ( .A(n343), .B(n344), .C(n345), .Z(n337) );
  GTECH_NOT U188 ( .A(n346), .Z(n342) );
  GTECH_XOR2 U189 ( .A(n346), .B(n347), .Z(n339) );
  GTECH_OAI21 U190 ( .A(b[14]), .B(a[14]), .C(n348), .Z(n346) );
  GTECH_OAI21 U191 ( .A(n349), .B(n345), .C(n350), .Z(sum[13]) );
  GTECH_MUX2 U192 ( .A(n351), .B(n352), .S(b[13]), .Z(n350) );
  GTECH_OR_NOT U193 ( .A(a[13]), .B(n349), .Z(n352) );
  GTECH_XOR2 U194 ( .A(a[13]), .B(n349), .Z(n351) );
  GTECH_OA21 U195 ( .A(n341), .B(n353), .C(n344), .Z(n349) );
  GTECH_OAI21 U196 ( .A(n341), .B(n354), .C(n355), .Z(sum[12]) );
  GTECH_AND_NOT U197 ( .A(n344), .B(n353), .Z(n354) );
  GTECH_NOT U198 ( .A(n356), .Z(n344) );
  GTECH_MUX2 U199 ( .A(n357), .B(n358), .S(n282), .Z(sum[11]) );
  GTECH_XOR2 U200 ( .A(n359), .B(n360), .Z(n358) );
  GTECH_XOR2 U201 ( .A(n361), .B(n362), .Z(n357) );
  GTECH_OA21 U202 ( .A(n363), .B(n364), .C(n365), .Z(n362) );
  GTECH_NOT U203 ( .A(n359), .Z(n361) );
  GTECH_XOR2 U204 ( .A(a[11]), .B(b[11]), .Z(n359) );
  GTECH_NOT U205 ( .A(n366), .Z(sum[10]) );
  GTECH_MUX2 U206 ( .A(n367), .B(n368), .S(n282), .Z(n366) );
  GTECH_XOR2 U207 ( .A(n369), .B(n370), .Z(n368) );
  GTECH_XOR2 U208 ( .A(n369), .B(n364), .Z(n367) );
  GTECH_OA21 U209 ( .A(n280), .B(n371), .C(n372), .Z(n364) );
  GTECH_OR_NOT U210 ( .A(n283), .B(b[8]), .Z(n371) );
  GTECH_AND_NOT U211 ( .A(n365), .B(n363), .Z(n369) );
  GTECH_XOR2 U212 ( .A(cin), .B(n306), .Z(sum[0]) );
  GTECH_NOT U213 ( .A(n373), .Z(n306) );
  GTECH_OAI21 U214 ( .A(n341), .B(n374), .C(n355), .Z(cout) );
  GTECH_OR3 U215 ( .A(n356), .B(n353), .C(n331), .Z(n355) );
  GTECH_NOT U216 ( .A(n341), .Z(n331) );
  GTECH_AND2 U217 ( .A(a[12]), .B(b[12]), .Z(n356) );
  GTECH_OA21 U218 ( .A(n333), .B(n338), .C(n375), .Z(n374) );
  GTECH_OAI21 U219 ( .A(a[15]), .B(n376), .C(b[15]), .Z(n375) );
  GTECH_NOT U220 ( .A(n333), .Z(n376) );
  GTECH_NOT U221 ( .A(a[15]), .Z(n338) );
  GTECH_OA21 U222 ( .A(n347), .B(n377), .C(n348), .Z(n333) );
  GTECH_NOT U223 ( .A(n336), .Z(n348) );
  GTECH_AND2 U224 ( .A(b[14]), .B(a[14]), .Z(n336) );
  GTECH_NOR2 U225 ( .A(b[14]), .B(a[14]), .Z(n377) );
  GTECH_OA21 U226 ( .A(n343), .B(n353), .C(n345), .Z(n347) );
  GTECH_OR_NOT U227 ( .A(n378), .B(b[13]), .Z(n345) );
  GTECH_NOR2 U228 ( .A(b[12]), .B(a[12]), .Z(n353) );
  GTECH_AND_NOT U229 ( .A(n378), .B(b[13]), .Z(n343) );
  GTECH_NOT U230 ( .A(a[13]), .Z(n378) );
  GTECH_AOI21 U231 ( .A(n282), .B(n379), .C(n286), .Z(n341) );
  GTECH_NOR2 U232 ( .A(n282), .B(n285), .Z(n286) );
  GTECH_XOR2 U233 ( .A(n280), .B(b[8]), .Z(n285) );
  GTECH_OA21 U234 ( .A(a[11]), .B(n360), .C(n380), .Z(n379) );
  GTECH_AO21 U235 ( .A(n360), .B(a[11]), .C(b[11]), .Z(n380) );
  GTECH_OAI21 U236 ( .A(n370), .B(n363), .C(n365), .Z(n360) );
  GTECH_OR_NOT U237 ( .A(n381), .B(a[10]), .Z(n365) );
  GTECH_NOT U238 ( .A(b[10]), .Z(n381) );
  GTECH_NOR2 U239 ( .A(b[10]), .B(a[10]), .Z(n363) );
  GTECH_OA21 U240 ( .A(n382), .B(n283), .C(n372), .Z(n370) );
  GTECH_NOT U241 ( .A(n284), .Z(n372) );
  GTECH_AND2 U242 ( .A(b[9]), .B(a[9]), .Z(n284) );
  GTECH_NOR2 U243 ( .A(b[9]), .B(a[9]), .Z(n283) );
  GTECH_AND2 U244 ( .A(n280), .B(n383), .Z(n382) );
  GTECH_NOT U245 ( .A(b[8]), .Z(n383) );
  GTECH_NOT U246 ( .A(a[8]), .Z(n280) );
  GTECH_MUX2 U247 ( .A(n311), .B(n384), .S(n289), .Z(n282) );
  GTECH_NOT U248 ( .A(n385), .Z(n289) );
  GTECH_MUX2 U249 ( .A(n386), .B(n373), .S(n307), .Z(n385) );
  GTECH_NOT U250 ( .A(cin), .Z(n307) );
  GTECH_XOR2 U251 ( .A(a[0]), .B(n328), .Z(n373) );
  GTECH_OA21 U252 ( .A(n308), .B(n309), .C(n310), .Z(n386) );
  GTECH_OAI21 U253 ( .A(a[3]), .B(n387), .C(b[3]), .Z(n310) );
  GTECH_NOT U254 ( .A(a[3]), .Z(n309) );
  GTECH_NOT U255 ( .A(n387), .Z(n308) );
  GTECH_ADD_ABC U256 ( .A(n322), .B(a[2]), .C(b[2]), .COUT(n387) );
  GTECH_AOI21 U257 ( .A(n388), .B(n327), .C(n389), .Z(n322) );
  GTECH_AOI21 U258 ( .A(n390), .B(a[1]), .C(b[1]), .Z(n389) );
  GTECH_NOT U259 ( .A(n327), .Z(n390) );
  GTECH_AND_NOT U260 ( .A(n328), .B(a[0]), .Z(n327) );
  GTECH_NOT U261 ( .A(b[0]), .Z(n328) );
  GTECH_NOT U262 ( .A(a[1]), .Z(n388) );
  GTECH_OA21 U263 ( .A(a[7]), .B(n291), .C(n391), .Z(n384) );
  GTECH_AO21 U264 ( .A(n291), .B(a[7]), .C(b[7]), .Z(n391) );
  GTECH_AO21 U265 ( .A(n298), .B(a[6]), .C(n392), .Z(n291) );
  GTECH_OA21 U266 ( .A(a[6]), .B(n298), .C(b[6]), .Z(n392) );
  GTECH_OAI21 U267 ( .A(n393), .B(n301), .C(n394), .Z(n298) );
  GTECH_NOT U268 ( .A(n300), .Z(n394) );
  GTECH_AND2 U269 ( .A(a[5]), .B(b[5]), .Z(n300) );
  GTECH_NOR2 U270 ( .A(a[5]), .B(b[5]), .Z(n301) );
  GTECH_NOR2 U271 ( .A(a[4]), .B(b[4]), .Z(n393) );
  GTECH_XOR2 U272 ( .A(a[4]), .B(b[4]), .Z(n311) );
endmodule

