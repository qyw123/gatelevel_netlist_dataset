
module frequency_counter ( clk, reset, signal, period, period_load, segments, 
        digit, dbg_state, dbg_clk_count, dbg_edge_count );
  input [11:0] period;
  output [6:0] segments;
  output [1:0] dbg_state;
  output [2:0] dbg_clk_count;
  output [2:0] dbg_edge_count;
  input clk, reset, signal, period_load;
  output digit;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21,
         update_digits, N62, N112, N114, N116, N118, N120, N122, N124, N126,
         N128, N130, N132, N133, N134, N136, N138, N140, N142, N144, N146,
         N147, N148, N150, N151, N152, N154, N156, N158, N159, N160, N162,
         N164, N166, N167, N168, N169, N170, edge_detect0_q2, edge_detect0_q1,
         edge_detect0_q0, seven_segment0_N22, seven_segment0_N20,
         seven_segment0_N18, seven_segment0_N16, seven_segment0_N14,
         seven_segment0_N12, seven_segment0_N10, seven_segment0_N9,
         seven_segment0_N8, seven_segment0_N6, n13, n14, n15, n16, n17, n21,
         n23, n26, n27, n28, n29, n31, n32, n33, n79, n160, sub_85_carry_2_,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334;
  wire   [8:0] clk_counter;
  wire   [3:0] edge_counter;
  wire   [11:0] update_period;
  wire   [3:0] ten_count;
  wire   [3:0] unit_count;
  wire   [0:3] seven_segment0_unit_count_reg;
  wire   [0:3] seven_segment0_ten_count_reg;

  GTECH_FJK1S update_period_reg_11_ ( .J(n79), .K(n79), .TI(N21), .TE(N20), 
        .CP(clk), .Q(update_period[11]) );
  GTECH_FJK1S update_period_reg_10_ ( .J(n79), .K(n79), .TI(N19), .TE(N20), 
        .CP(clk), .Q(update_period[10]) );
  GTECH_FJK1S update_period_reg_9_ ( .J(n79), .K(n79), .TI(N18), .TE(N20), 
        .CP(clk), .Q(update_period[9]) );
  GTECH_FJK1S update_period_reg_8_ ( .J(n79), .K(n79), .TI(N17), .TE(N20), 
        .CP(clk), .Q(update_period[8]) );
  GTECH_FJK1S update_period_reg_7_ ( .J(n79), .K(n79), .TI(N16), .TE(N20), 
        .CP(clk), .Q(update_period[7]) );
  GTECH_FJK1S update_period_reg_6_ ( .J(n79), .K(n79), .TI(N15), .TE(N20), 
        .CP(clk), .Q(update_period[6]) );
  GTECH_FJK1S update_period_reg_5_ ( .J(n79), .K(n79), .TI(N14), .TE(N20), 
        .CP(clk), .Q(update_period[5]) );
  GTECH_FJK1S update_period_reg_4_ ( .J(n79), .K(n79), .TI(N13), .TE(N20), 
        .CP(clk), .Q(update_period[4]) );
  GTECH_FJK1S update_period_reg_3_ ( .J(n79), .K(n79), .TI(N12), .TE(N20), 
        .CP(clk), .Q(update_period[3]) );
  GTECH_FJK1S update_period_reg_2_ ( .J(n79), .K(n79), .TI(N11), .TE(N20), 
        .CP(clk), .Q(update_period[2]) );
  GTECH_FJK1S update_period_reg_1_ ( .J(n79), .K(n79), .TI(N10), .TE(N20), 
        .CP(clk), .Q(update_period[1]) );
  GTECH_FJK1S update_period_reg_0_ ( .J(n79), .K(n79), .TI(N9), .TE(N20), .CP(
        clk), .Q(update_period[0]), .QN(n176) );
  GTECH_FD1 edge_detect0_q0_reg ( .D(signal), .CP(clk), .Q(edge_detect0_q0) );
  GTECH_FD1 edge_detect0_q1_reg ( .D(edge_detect0_q0), .CP(clk), .Q(
        edge_detect0_q1) );
  GTECH_FD1 edge_detect0_q2_reg ( .D(edge_detect0_q1), .CP(clk), .Q(
        edge_detect0_q2), .QN(n13) );
  GTECH_FJK1S edge_counter_reg_5_ ( .J(n79), .K(n79), .TI(N146), .TE(N147), 
        .CP(clk), .Q(dbg_edge_count[1]), .QN(n175) );
  GTECH_FJK1S edge_counter_reg_6_ ( .J(n79), .K(n79), .TI(N148), .TE(N147), 
        .CP(clk), .Q(dbg_edge_count[2]), .QN(n174) );
  GTECH_FJK1S state_reg_0_ ( .J(n79), .K(n79), .TI(N150), .TE(N151), .CP(clk), 
        .Q(dbg_state[0]), .QN(n14) );
  GTECH_FJK1S state_reg_1_ ( .J(n79), .K(n79), .TI(N152), .TE(N151), .CP(clk), 
        .Q(dbg_state[1]), .QN(n15) );
  GTECH_FJK1S clk_counter_reg_10_ ( .J(n79), .K(n79), .TI(N132), .TE(N133), 
        .CP(clk), .Q(dbg_clk_count[1]), .QN(n173) );
  GTECH_FJK1S clk_counter_reg_0_ ( .J(n79), .K(n79), .TI(N112), .TE(N133), 
        .CP(clk), .Q(clk_counter[0]), .QN(n172) );
  GTECH_FJK1S clk_counter_reg_1_ ( .J(n79), .K(n79), .TI(N114), .TE(N133), 
        .CP(clk), .Q(clk_counter[1]), .QN(n171) );
  GTECH_FJK1S clk_counter_reg_2_ ( .J(n79), .K(n79), .TI(N116), .TE(N133), 
        .CP(clk), .Q(clk_counter[2]), .QN(n170) );
  GTECH_FJK1S clk_counter_reg_3_ ( .J(n79), .K(n79), .TI(N118), .TE(N133), 
        .CP(clk), .Q(clk_counter[3]), .QN(n169) );
  GTECH_FJK1S clk_counter_reg_4_ ( .J(n79), .K(n79), .TI(N120), .TE(N133), 
        .CP(clk), .Q(clk_counter[4]), .QN(n168) );
  GTECH_FJK1S clk_counter_reg_5_ ( .J(n79), .K(n79), .TI(N122), .TE(N133), 
        .CP(clk), .Q(clk_counter[5]), .QN(n167) );
  GTECH_FJK1S clk_counter_reg_6_ ( .J(n79), .K(n79), .TI(N124), .TE(N133), 
        .CP(clk), .Q(clk_counter[6]), .QN(n166) );
  GTECH_FJK1S clk_counter_reg_7_ ( .J(n79), .K(n79), .TI(N126), .TE(N133), 
        .CP(clk), .Q(clk_counter[7]), .QN(n165) );
  GTECH_FJK1S clk_counter_reg_8_ ( .J(n79), .K(n79), .TI(N128), .TE(N133), 
        .CP(clk), .Q(clk_counter[8]), .QN(n164) );
  GTECH_FJK1S clk_counter_reg_9_ ( .J(n79), .K(n79), .TI(N130), .TE(N133), 
        .CP(clk), .Q(dbg_clk_count[0]), .QN(n163) );
  GTECH_FJK1S clk_counter_reg_11_ ( .J(n79), .K(n79), .TI(N134), .TE(N133), 
        .CP(clk), .Q(dbg_clk_count[2]), .QN(n162) );
  GTECH_FJK1S update_digits_reg ( .J(n79), .K(n79), .TI(N170), .TE(N169), .CP(
        clk), .Q(update_digits), .QN(n16) );
  GTECH_FJK1S edge_counter_reg_4_ ( .J(n79), .K(n79), .TI(N144), .TE(N147), 
        .CP(clk), .Q(dbg_edge_count[0]), .QN(n161) );
  GTECH_FJK1S edge_counter_reg_0_ ( .J(n79), .K(n79), .TI(N136), .TE(N147), 
        .CP(clk), .Q(N62), .QN(n17) );
  GTECH_FJK1S unit_count_reg_0_ ( .J(n79), .K(n79), .TI(N162), .TE(N167), .CP(
        clk), .Q(unit_count[0]) );
  GTECH_FJK1S edge_counter_reg_1_ ( .J(n79), .K(n79), .TI(N138), .TE(N147), 
        .CP(clk), .Q(sub_85_carry_2_) );
  GTECH_FJK1S unit_count_reg_1_ ( .J(n79), .K(n79), .TI(N164), .TE(N167), .CP(
        clk), .Q(unit_count[1]) );
  GTECH_FJK1S edge_counter_reg_2_ ( .J(n79), .K(n79), .TI(N140), .TE(N147), 
        .CP(clk), .Q(edge_counter[2]), .QN(n21) );
  GTECH_FJK1S unit_count_reg_2_ ( .J(n79), .K(n79), .TI(N166), .TE(N167), .CP(
        clk), .Q(unit_count[2]) );
  GTECH_FJK1S edge_counter_reg_3_ ( .J(n79), .K(n79), .TI(N142), .TE(N147), 
        .CP(clk), .Q(edge_counter[3]), .QN(n23) );
  GTECH_FJK1S unit_count_reg_3_ ( .J(n79), .K(n79), .TI(N168), .TE(N167), .CP(
        clk), .Q(unit_count[3]) );
  GTECH_FJK1S ten_count_reg_0_ ( .J(n79), .K(n79), .TI(N154), .TE(N159), .CP(
        clk), .Q(ten_count[0]) );
  GTECH_FJK1S ten_count_reg_1_ ( .J(n79), .K(n79), .TI(N156), .TE(N159), .CP(
        clk), .Q(ten_count[1]) );
  GTECH_FJK1S ten_count_reg_2_ ( .J(n79), .K(n79), .TI(N158), .TE(N159), .CP(
        clk), .Q(ten_count[2]) );
  GTECH_FJK1S ten_count_reg_3_ ( .J(n79), .K(n79), .TI(N160), .TE(N159), .CP(
        clk), .Q(n26) );
  GTECH_FJK1S seven_segment0_unit_count_reg_reg_0_ ( .J(n79), .K(n79), .TI(
        seven_segment0_N16), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_unit_count_reg[0]), .QN(n27) );
  GTECH_FJK1S seven_segment0_unit_count_reg_reg_1_ ( .J(n79), .K(n79), .TI(
        seven_segment0_N18), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_unit_count_reg[1]), .QN(n28) );
  GTECH_FJK1S seven_segment0_unit_count_reg_reg_2_ ( .J(n79), .K(n79), .TI(
        seven_segment0_N20), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_unit_count_reg[2]), .QN(n29) );
  GTECH_FJK1S seven_segment0_unit_count_reg_reg_3_ ( .J(n79), .K(n79), .TI(
        seven_segment0_N22), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_unit_count_reg[3]) );
  GTECH_FJK1S seven_segment0_ten_count_reg_reg_0_ ( .J(n79), .K(n79), .TI(
        seven_segment0_N8), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_ten_count_reg[0]), .QN(n31) );
  GTECH_FJK1S seven_segment0_ten_count_reg_reg_1_ ( .J(n79), .K(n79), .TI(
        seven_segment0_N10), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_ten_count_reg[1]), .QN(n32) );
  GTECH_FJK1S seven_segment0_ten_count_reg_reg_2_ ( .J(n79), .K(n79), .TI(
        seven_segment0_N12), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_ten_count_reg[2]), .QN(n33) );
  GTECH_FJK1S seven_segment0_ten_count_reg_reg_3_ ( .J(n79), .K(n79), .TI(
        seven_segment0_N14), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_ten_count_reg[3]) );
  GTECH_FD1 seven_segment0_digit_reg ( .D(seven_segment0_N6), .CP(clk), .Q(
        digit), .QN(n160) );
  GTECH_ZERO U168 ( .Z(n79) );
  GTECH_OR_NOT U169 ( .A(reset), .B(n16), .Z(seven_segment0_N9) );
  GTECH_AND2 U170 ( .A(ten_count[0]), .B(n188), .Z(seven_segment0_N8) );
  GTECH_AND2 U171 ( .A(n160), .B(n188), .Z(seven_segment0_N6) );
  GTECH_AND2 U172 ( .A(unit_count[3]), .B(n188), .Z(seven_segment0_N22) );
  GTECH_AND2 U173 ( .A(unit_count[2]), .B(n188), .Z(seven_segment0_N20) );
  GTECH_AND2 U174 ( .A(unit_count[1]), .B(n188), .Z(seven_segment0_N18) );
  GTECH_AND2 U175 ( .A(unit_count[0]), .B(n188), .Z(seven_segment0_N16) );
  GTECH_AND2 U176 ( .A(n26), .B(n188), .Z(seven_segment0_N14) );
  GTECH_AND2 U177 ( .A(ten_count[2]), .B(n188), .Z(seven_segment0_N12) );
  GTECH_AND2 U178 ( .A(ten_count[1]), .B(n188), .Z(seven_segment0_N10) );
  GTECH_OR_NOT U179 ( .A(n189), .B(n190), .Z(segments[6]) );
  GTECH_NOT U180 ( .A(n191), .Z(n189) );
  GTECH_OR_NOT U181 ( .A(n192), .B(n190), .Z(segments[5]) );
  GTECH_NOT U182 ( .A(n193), .Z(n190) );
  GTECH_OAI21 U183 ( .A(n194), .B(n195), .C(n196), .Z(n193) );
  GTECH_NOT U184 ( .A(n197), .Z(n192) );
  GTECH_NAND3 U185 ( .A(n191), .B(n198), .C(n199), .Z(segments[3]) );
  GTECH_NOT U186 ( .A(segments[4]), .Z(n198) );
  GTECH_OAI21 U187 ( .A(n200), .B(n201), .C(n197), .Z(segments[4]) );
  GTECH_NAND3 U188 ( .A(n196), .B(n195), .C(n202), .Z(segments[2]) );
  GTECH_AND3 U189 ( .A(n203), .B(n204), .C(n199), .Z(n196) );
  GTECH_NAND3 U190 ( .A(n205), .B(n206), .C(n207), .Z(n204) );
  GTECH_NAND3 U191 ( .A(n203), .B(n191), .C(n208), .Z(segments[1]) );
  GTECH_OA21 U192 ( .A(n206), .B(n200), .C(n195), .Z(n208) );
  GTECH_NAND4 U193 ( .A(n206), .B(n209), .C(n205), .D(n194), .Z(n203) );
  GTECH_NAND3 U194 ( .A(n199), .B(n191), .C(n210), .Z(segments[0]) );
  GTECH_OA21 U195 ( .A(n194), .B(n195), .C(n202), .Z(n210) );
  GTECH_NOT U196 ( .A(n211), .Z(n202) );
  GTECH_OAI21 U197 ( .A(n206), .B(n200), .C(n197), .Z(n211) );
  GTECH_OR_NOT U198 ( .A(n201), .B(n212), .Z(n197) );
  GTECH_NOT U199 ( .A(n195), .Z(n212) );
  GTECH_OR_NOT U200 ( .A(n205), .B(n209), .Z(n195) );
  GTECH_OR_NOT U201 ( .A(n205), .B(n207), .Z(n191) );
  GTECH_NOT U202 ( .A(n200), .Z(n207) );
  GTECH_OR_NOT U203 ( .A(n213), .B(n214), .Z(n200) );
  GTECH_NOT U204 ( .A(n209), .Z(n214) );
  GTECH_NAND4 U205 ( .A(n209), .B(n201), .C(n205), .D(n194), .Z(n199) );
  GTECH_NOT U206 ( .A(n213), .Z(n194) );
  GTECH_MUX2 U207 ( .A(seven_segment0_ten_count_reg[3]), .B(
        seven_segment0_unit_count_reg[3]), .S(n160), .Z(n213) );
  GTECH_NOT U208 ( .A(n215), .Z(n205) );
  GTECH_MUX2 U209 ( .A(n33), .B(n29), .S(n160), .Z(n215) );
  GTECH_NOT U210 ( .A(n206), .Z(n201) );
  GTECH_MUX2 U211 ( .A(n31), .B(n27), .S(n160), .Z(n206) );
  GTECH_MUX2 U212 ( .A(n32), .B(n28), .S(n160), .Z(n209) );
  GTECH_AO21 U213 ( .A(period[0]), .B(n216), .C(reset), .Z(N9) );
  GTECH_AND2 U214 ( .A(period[11]), .B(n216), .Z(N21) );
  GTECH_OR_NOT U215 ( .A(n216), .B(n188), .Z(N20) );
  GTECH_AO21 U216 ( .A(period[10]), .B(n216), .C(reset), .Z(N19) );
  GTECH_AND2 U217 ( .A(period[9]), .B(n216), .Z(N18) );
  GTECH_AND2 U218 ( .A(period[8]), .B(n216), .Z(N17) );
  GTECH_AND2 U219 ( .A(N170), .B(n217), .Z(N168) );
  GTECH_OR_NOT U220 ( .A(n218), .B(n219), .Z(N167) );
  GTECH_AND2 U221 ( .A(N170), .B(n220), .Z(N166) );
  GTECH_AND2 U222 ( .A(sub_85_carry_2_), .B(N170), .Z(N164) );
  GTECH_AND2 U223 ( .A(N170), .B(n221), .Z(N162) );
  GTECH_NOT U224 ( .A(n222), .Z(N170) );
  GTECH_OR_NOT U225 ( .A(reset), .B(n218), .Z(n222) );
  GTECH_NOT U226 ( .A(n223), .Z(n218) );
  GTECH_MUX2 U227 ( .A(n224), .B(n225), .S(n26), .Z(N160) );
  GTECH_OAI21 U228 ( .A(ten_count[2]), .B(n226), .C(n227), .Z(n225) );
  GTECH_NOT U229 ( .A(n228), .Z(n227) );
  GTECH_AND2 U230 ( .A(n229), .B(ten_count[2]), .Z(n224) );
  GTECH_AO21 U231 ( .A(period[7]), .B(n216), .C(reset), .Z(N16) );
  GTECH_OAI21 U232 ( .A(n230), .B(n231), .C(n232), .Z(N159) );
  GTECH_MUX2 U233 ( .A(n229), .B(n228), .S(ten_count[2]), .Z(N158) );
  GTECH_OAI21 U234 ( .A(ten_count[1]), .B(n226), .C(n233), .Z(n228) );
  GTECH_NOT U235 ( .A(n234), .Z(n229) );
  GTECH_NAND3 U236 ( .A(ten_count[1]), .B(ten_count[0]), .C(N152), .Z(n234) );
  GTECH_MUX2 U237 ( .A(n235), .B(N154), .S(ten_count[1]), .Z(N156) );
  GTECH_AND2 U238 ( .A(N152), .B(ten_count[0]), .Z(n235) );
  GTECH_NOT U239 ( .A(n233), .Z(N154) );
  GTECH_OR_NOT U240 ( .A(ten_count[0]), .B(N152), .Z(n233) );
  GTECH_OR_NOT U241 ( .A(n236), .B(n237), .Z(N151) );
  GTECH_OA21 U242 ( .A(n14), .B(n238), .C(n219), .Z(n237) );
  GTECH_NOT U243 ( .A(n239), .Z(n219) );
  GTECH_OAI21 U244 ( .A(n240), .B(n230), .C(n188), .Z(n239) );
  GTECH_AND2 U245 ( .A(period[6]), .B(n216), .Z(N15) );
  GTECH_OAI21 U246 ( .A(n226), .B(n238), .C(n241), .Z(N148) );
  GTECH_MUX2 U247 ( .A(n242), .B(n243), .S(n174), .Z(n241) );
  GTECH_OR3 U248 ( .A(n175), .B(n244), .C(n245), .Z(n243) );
  GTECH_AND_NOT U249 ( .A(n246), .B(n247), .Z(n242) );
  GTECH_MUX2 U250 ( .A(n226), .B(n244), .S(n175), .Z(n246) );
  GTECH_NAND3 U251 ( .A(n248), .B(n223), .C(n232), .Z(N147) );
  GTECH_OA21 U252 ( .A(n236), .B(n249), .C(n188), .Z(n232) );
  GTECH_OR_NOT U253 ( .A(n14), .B(n238), .Z(n249) );
  GTECH_NAND4 U254 ( .A(n175), .B(n174), .C(n161), .D(n250), .Z(n238) );
  GTECH_NOT U255 ( .A(n15), .Z(n236) );
  GTECH_OR_NOT U256 ( .A(n15), .B(n14), .Z(n223) );
  GTECH_NAND3 U257 ( .A(n14), .B(edge_detect0_q1), .C(n13), .Z(n248) );
  GTECH_MUX2 U258 ( .A(n247), .B(n251), .S(n175), .Z(N146) );
  GTECH_OAI21 U259 ( .A(n245), .B(n244), .C(n252), .Z(n251) );
  GTECH_OAI21 U260 ( .A(n253), .B(n244), .C(n254), .Z(n247) );
  GTECH_AO21 U261 ( .A(n250), .B(n161), .C(n226), .Z(n254) );
  GTECH_NOT U262 ( .A(n245), .Z(n253) );
  GTECH_NAND3 U263 ( .A(n255), .B(n217), .C(n256), .Z(n245) );
  GTECH_NOT U264 ( .A(n161), .Z(n255) );
  GTECH_OR_NOT U265 ( .A(n257), .B(n252), .Z(N144) );
  GTECH_NAND3 U266 ( .A(N152), .B(n250), .C(n161), .Z(n252) );
  GTECH_MUX2 U267 ( .A(n258), .B(n259), .S(n161), .Z(n257) );
  GTECH_AND3 U268 ( .A(n217), .B(N150), .C(n256), .Z(n259) );
  GTECH_NOT U269 ( .A(n23), .Z(n217) );
  GTECH_OAI21 U270 ( .A(n250), .B(n226), .C(n260), .Z(n258) );
  GTECH_OAI21 U271 ( .A(n23), .B(n261), .C(N150), .Z(n260) );
  GTECH_OR_NOT U272 ( .A(n23), .B(n262), .Z(n250) );
  GTECH_OAI21 U273 ( .A(n244), .B(n263), .C(n264), .Z(N142) );
  GTECH_MUX2 U274 ( .A(n265), .B(n266), .S(n23), .Z(n264) );
  GTECH_OR_NOT U275 ( .A(n267), .B(N152), .Z(n266) );
  GTECH_NOT U276 ( .A(n226), .Z(N152) );
  GTECH_XOR2 U277 ( .A(n23), .B(n256), .Z(n263) );
  GTECH_NOT U278 ( .A(n261), .Z(n256) );
  GTECH_NAND3 U279 ( .A(n221), .B(n220), .C(sub_85_carry_2_), .Z(n261) );
  GTECH_NOT U280 ( .A(n21), .Z(n220) );
  GTECH_OR_NOT U281 ( .A(n268), .B(n269), .Z(N140) );
  GTECH_MUX2 U282 ( .A(n270), .B(n271), .S(n21), .Z(n269) );
  GTECH_NAND3 U283 ( .A(sub_85_carry_2_), .B(n221), .C(N150), .Z(n271) );
  GTECH_NOT U284 ( .A(n244), .Z(N150) );
  GTECH_NOT U285 ( .A(n17), .Z(n221) );
  GTECH_AND2 U286 ( .A(n272), .B(n273), .Z(n270) );
  GTECH_MUX2 U287 ( .A(n244), .B(n226), .S(sub_85_carry_2_), .Z(n272) );
  GTECH_NOT U288 ( .A(n265), .Z(n268) );
  GTECH_OR_NOT U289 ( .A(n226), .B(n267), .Z(n265) );
  GTECH_NOT U290 ( .A(n262), .Z(n267) );
  GTECH_OR_NOT U291 ( .A(sub_85_carry_2_), .B(n21), .Z(n262) );
  GTECH_AO21 U292 ( .A(period[5]), .B(n216), .C(reset), .Z(N14) );
  GTECH_MUX2 U293 ( .A(n274), .B(n275), .S(sub_85_carry_2_), .Z(N138) );
  GTECH_NOT U294 ( .A(n273), .Z(n275) );
  GTECH_OAI21 U295 ( .A(n17), .B(n244), .C(n226), .Z(n274) );
  GTECH_OAI21 U296 ( .A(n17), .B(n226), .C(n273), .Z(N136) );
  GTECH_OR_NOT U297 ( .A(n244), .B(n17), .Z(n273) );
  GTECH_OR_NOT U298 ( .A(reset), .B(n276), .Z(n244) );
  GTECH_OR_NOT U299 ( .A(N169), .B(n15), .Z(n226) );
  GTECH_OR_NOT U300 ( .A(n14), .B(n188), .Z(N169) );
  GTECH_AND2 U301 ( .A(n277), .B(n278), .Z(N134) );
  GTECH_OAI21 U302 ( .A(n173), .B(n279), .C(n162), .Z(n278) );
  GTECH_OR_NOT U303 ( .A(n276), .B(n188), .Z(N133) );
  GTECH_NOT U304 ( .A(reset), .Z(n188) );
  GTECH_NOT U305 ( .A(n231), .Z(n276) );
  GTECH_OR_NOT U306 ( .A(n240), .B(n15), .Z(n231) );
  GTECH_NOT U307 ( .A(n14), .Z(n240) );
  GTECH_AND2 U308 ( .A(n280), .B(n277), .Z(N132) );
  GTECH_XOR2 U309 ( .A(n279), .B(n173), .Z(n280) );
  GTECH_OR_NOT U310 ( .A(n163), .B(n281), .Z(n279) );
  GTECH_NOT U311 ( .A(n282), .Z(n281) );
  GTECH_AND2 U312 ( .A(n283), .B(n277), .Z(N130) );
  GTECH_XOR2 U313 ( .A(n282), .B(n163), .Z(n283) );
  GTECH_OR_NOT U314 ( .A(n164), .B(n284), .Z(n282) );
  GTECH_NOT U315 ( .A(n285), .Z(n284) );
  GTECH_AND2 U316 ( .A(period[4]), .B(n216), .Z(N13) );
  GTECH_AND2 U317 ( .A(n286), .B(n277), .Z(N128) );
  GTECH_XOR2 U318 ( .A(n285), .B(n164), .Z(n286) );
  GTECH_OR_NOT U319 ( .A(n165), .B(n287), .Z(n285) );
  GTECH_NOT U320 ( .A(n288), .Z(n287) );
  GTECH_AND2 U321 ( .A(n289), .B(n277), .Z(N126) );
  GTECH_XOR2 U322 ( .A(n288), .B(n165), .Z(n289) );
  GTECH_OR_NOT U323 ( .A(n166), .B(n290), .Z(n288) );
  GTECH_NOT U324 ( .A(n291), .Z(n290) );
  GTECH_AND2 U325 ( .A(n292), .B(n277), .Z(N124) );
  GTECH_XOR2 U326 ( .A(n291), .B(n166), .Z(n292) );
  GTECH_OR_NOT U327 ( .A(n167), .B(n293), .Z(n291) );
  GTECH_NOT U328 ( .A(n294), .Z(n293) );
  GTECH_AND2 U329 ( .A(n295), .B(n277), .Z(N122) );
  GTECH_XOR2 U330 ( .A(n294), .B(n167), .Z(n295) );
  GTECH_OR_NOT U331 ( .A(n168), .B(n296), .Z(n294) );
  GTECH_NOT U332 ( .A(n297), .Z(n296) );
  GTECH_AND2 U333 ( .A(n298), .B(n277), .Z(N120) );
  GTECH_XOR2 U334 ( .A(n297), .B(n168), .Z(n298) );
  GTECH_OR_NOT U335 ( .A(n169), .B(n299), .Z(n297) );
  GTECH_NOT U336 ( .A(n300), .Z(n299) );
  GTECH_AO21 U337 ( .A(period[3]), .B(n216), .C(reset), .Z(N12) );
  GTECH_AND2 U338 ( .A(n301), .B(n277), .Z(N118) );
  GTECH_XOR2 U339 ( .A(n300), .B(n169), .Z(n301) );
  GTECH_NAND3 U340 ( .A(n302), .B(n303), .C(n304), .Z(n300) );
  GTECH_NOT U341 ( .A(n170), .Z(n304) );
  GTECH_OAI22 U342 ( .A(n170), .B(n305), .C(n306), .D(n307), .Z(N116) );
  GTECH_MUX2 U343 ( .A(n302), .B(n308), .S(n170), .Z(n307) );
  GTECH_OR_NOT U344 ( .A(n172), .B(n302), .Z(n308) );
  GTECH_MUX2 U345 ( .A(N112), .B(n309), .S(n171), .Z(N114) );
  GTECH_AND2 U346 ( .A(n277), .B(n303), .Z(n309) );
  GTECH_NOT U347 ( .A(n305), .Z(N112) );
  GTECH_OR_NOT U348 ( .A(n303), .B(n277), .Z(n305) );
  GTECH_NOT U349 ( .A(n306), .Z(n277) );
  GTECH_OR_NOT U350 ( .A(reset), .B(n230), .Z(n306) );
  GTECH_OAI21 U351 ( .A(n310), .B(n311), .C(n312), .Z(n230) );
  GTECH_AOI2N2 U352 ( .A(update_period[11]), .B(n162), .C(n313), .D(n314), .Z(
        n312) );
  GTECH_AOI222 U353 ( .A(update_period[9]), .B(n163), .C(n315), .D(
        update_period[8]), .E(update_period[10]), .F(n173), .Z(n314) );
  GTECH_OA21 U354 ( .A(n163), .B(update_period[9]), .C(n164), .Z(n315) );
  GTECH_OAI21 U355 ( .A(update_period[8]), .B(n164), .C(n316), .Z(n311) );
  GTECH_NOT U356 ( .A(n313), .Z(n316) );
  GTECH_OAI22 U357 ( .A(update_period[10]), .B(n173), .C(update_period[11]), 
        .D(n162), .Z(n313) );
  GTECH_OAI22 U358 ( .A(update_period[9]), .B(n163), .C(n317), .D(n318), .Z(
        n310) );
  GTECH_OAI22 U359 ( .A(n319), .B(n320), .C(n321), .D(n319), .Z(n318) );
  GTECH_AOI22 U360 ( .A(n168), .B(update_period[4]), .C(update_period[5]), .D(
        n167), .Z(n321) );
  GTECH_OAI22 U361 ( .A(update_period[4]), .B(n168), .C(n322), .D(n323), .Z(
        n320) );
  GTECH_AO22 U362 ( .A(n324), .B(n170), .C(n169), .D(update_period[3]), .Z(
        n323) );
  GTECH_AND2 U363 ( .A(n325), .B(update_period[2]), .Z(n324) );
  GTECH_AND3 U364 ( .A(n326), .B(n327), .C(n325), .Z(n322) );
  GTECH_OR_NOT U365 ( .A(n169), .B(n328), .Z(n325) );
  GTECH_NOT U366 ( .A(update_period[3]), .Z(n328) );
  GTECH_OAI22 U367 ( .A(n302), .B(n329), .C(n303), .D(n176), .Z(n327) );
  GTECH_AOI2N2 U368 ( .A(n302), .B(n329), .C(n170), .D(update_period[2]), .Z(
        n326) );
  GTECH_NOT U369 ( .A(update_period[1]), .Z(n329) );
  GTECH_NOT U370 ( .A(n171), .Z(n302) );
  GTECH_OAI21 U371 ( .A(update_period[5]), .B(n167), .C(n330), .Z(n319) );
  GTECH_OA21 U372 ( .A(update_period[6]), .B(n166), .C(n331), .Z(n330) );
  GTECH_AO22 U373 ( .A(n332), .B(n166), .C(n165), .D(update_period[7]), .Z(
        n317) );
  GTECH_AND2 U374 ( .A(n331), .B(update_period[6]), .Z(n332) );
  GTECH_OR_NOT U375 ( .A(n165), .B(n333), .Z(n331) );
  GTECH_NOT U376 ( .A(update_period[7]), .Z(n333) );
  GTECH_NOT U377 ( .A(n172), .Z(n303) );
  GTECH_AO21 U378 ( .A(period[2]), .B(n216), .C(reset), .Z(N11) );
  GTECH_AO21 U379 ( .A(period[1]), .B(n216), .C(reset), .Z(N10) );
  GTECH_NOT U380 ( .A(n334), .Z(n216) );
  GTECH_OR_NOT U381 ( .A(reset), .B(period_load), .Z(n334) );
endmodule

