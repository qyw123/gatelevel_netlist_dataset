
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_OR_NOT U83 ( .A(n97), .B(n93), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n98), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n98) );
  GTECH_OAI21 U86 ( .A(n99), .B(n100), .C(n101), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  GTECH_NOT U88 ( .A(n103), .Z(n99) );
  GTECH_OR_NOT U89 ( .A(n105), .B(I_b[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n106), .Z(n84) );
  GTECH_OR_NOT U91 ( .A(n107), .B(n108), .Z(n106) );
  GTECH_XOR2 U92 ( .A(n109), .B(n108), .Z(N153) );
  GTECH_NOT U93 ( .A(n110), .Z(n108) );
  GTECH_XOR3 U94 ( .A(n97), .B(n93), .C(n95), .Z(n110) );
  GTECH_XOR3 U95 ( .A(n102), .B(n104), .C(n103), .Z(n95) );
  GTECH_OAI21 U96 ( .A(n111), .B(n112), .C(n113), .Z(n103) );
  GTECH_OAI21 U97 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_NOT U98 ( .A(n115), .Z(n111) );
  GTECH_NOT U99 ( .A(n117), .Z(n104) );
  GTECH_OR_NOT U100 ( .A(n118), .B(I_b[7]), .Z(n117) );
  GTECH_NOT U101 ( .A(n100), .Z(n102) );
  GTECH_OR_NOT U102 ( .A(n119), .B(I_a[7]), .Z(n100) );
  GTECH_NOT U103 ( .A(I_b[6]), .Z(n119) );
  GTECH_ADD_ABC U104 ( .A(n120), .B(n121), .C(n122), .COUT(n93) );
  GTECH_NOT U105 ( .A(n123), .Z(n122) );
  GTECH_XOR2 U106 ( .A(n124), .B(n125), .Z(n121) );
  GTECH_AND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n125) );
  GTECH_NOT U108 ( .A(n94), .Z(n97) );
  GTECH_OR_NOT U109 ( .A(n124), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U110 ( .A(n107), .Z(n109) );
  GTECH_OR_NOT U111 ( .A(n126), .B(n127), .Z(n107) );
  GTECH_XOR2 U112 ( .A(n126), .B(n128), .Z(N152) );
  GTECH_NOT U113 ( .A(n127), .Z(n128) );
  GTECH_XNOR4 U114 ( .A(n124), .B(n123), .C(n129), .D(n120), .Z(n127) );
  GTECH_ADD_ABC U115 ( .A(n130), .B(n131), .C(n132), .COUT(n120) );
  GTECH_NOT U116 ( .A(n133), .Z(n132) );
  GTECH_XOR3 U117 ( .A(n134), .B(n135), .C(n136), .Z(n131) );
  GTECH_OR_NOT U118 ( .A(n137), .B(I_a[7]), .Z(n129) );
  GTECH_XOR3 U119 ( .A(n114), .B(n116), .C(n115), .Z(n123) );
  GTECH_OAI21 U120 ( .A(n138), .B(n139), .C(n140), .Z(n115) );
  GTECH_OAI21 U121 ( .A(n141), .B(n142), .C(n143), .Z(n140) );
  GTECH_NOT U122 ( .A(n142), .Z(n138) );
  GTECH_NOT U123 ( .A(n144), .Z(n116) );
  GTECH_OR_NOT U124 ( .A(n145), .B(I_b[7]), .Z(n144) );
  GTECH_NOT U125 ( .A(n112), .Z(n114) );
  GTECH_OR_NOT U126 ( .A(n118), .B(I_b[6]), .Z(n112) );
  GTECH_NOT U127 ( .A(I_a[6]), .Z(n118) );
  GTECH_OA21 U128 ( .A(n136), .B(n146), .C(n147), .Z(n124) );
  GTECH_OAI21 U129 ( .A(n134), .B(n148), .C(n135), .Z(n147) );
  GTECH_NOT U130 ( .A(n148), .Z(n136) );
  GTECH_ADD_ABC U131 ( .A(n149), .B(n150), .C(n151), .COUT(n126) );
  GTECH_NOT U132 ( .A(n152), .Z(n151) );
  GTECH_OA22 U133 ( .A(n153), .B(n105), .C(n154), .D(n155), .Z(n150) );
  GTECH_OA21 U134 ( .A(n156), .B(n157), .C(n158), .Z(n149) );
  GTECH_XOR3 U135 ( .A(n159), .B(n152), .C(n160), .Z(N151) );
  GTECH_OA21 U136 ( .A(n156), .B(n157), .C(n158), .Z(n160) );
  GTECH_OAI21 U137 ( .A(n161), .B(n162), .C(n163), .Z(n158) );
  GTECH_XOR2 U138 ( .A(n164), .B(n130), .Z(n152) );
  GTECH_ADD_ABC U139 ( .A(n165), .B(n166), .C(n167), .COUT(n130) );
  GTECH_NOT U140 ( .A(n168), .Z(n167) );
  GTECH_XOR3 U141 ( .A(n169), .B(n170), .C(n171), .Z(n166) );
  GTECH_XNOR4 U142 ( .A(n135), .B(n148), .C(n133), .D(n134), .Z(n164) );
  GTECH_NOT U143 ( .A(n146), .Z(n134) );
  GTECH_OR_NOT U144 ( .A(n172), .B(I_a[7]), .Z(n146) );
  GTECH_XOR3 U145 ( .A(n141), .B(n143), .C(n142), .Z(n133) );
  GTECH_OAI21 U146 ( .A(n173), .B(n174), .C(n175), .Z(n142) );
  GTECH_OAI21 U147 ( .A(n176), .B(n177), .C(n178), .Z(n175) );
  GTECH_NOT U148 ( .A(n177), .Z(n173) );
  GTECH_NOT U149 ( .A(n179), .Z(n143) );
  GTECH_OR_NOT U150 ( .A(n180), .B(I_b[7]), .Z(n179) );
  GTECH_NOT U151 ( .A(n139), .Z(n141) );
  GTECH_OR_NOT U152 ( .A(n145), .B(I_b[6]), .Z(n139) );
  GTECH_NOT U153 ( .A(I_a[5]), .Z(n145) );
  GTECH_OAI21 U154 ( .A(n171), .B(n181), .C(n182), .Z(n148) );
  GTECH_OAI21 U155 ( .A(n169), .B(n183), .C(n170), .Z(n182) );
  GTECH_NOT U156 ( .A(n183), .Z(n171) );
  GTECH_NOT U157 ( .A(n184), .Z(n135) );
  GTECH_OR_NOT U158 ( .A(n137), .B(I_a[6]), .Z(n184) );
  GTECH_OA22 U159 ( .A(n153), .B(n105), .C(n154), .D(n155), .Z(n159) );
  GTECH_NOT U160 ( .A(n185), .Z(n155) );
  GTECH_NOT U161 ( .A(I_a[7]), .Z(n105) );
  GTECH_XOR3 U162 ( .A(n156), .B(n161), .C(n186), .Z(N150) );
  GTECH_NOT U163 ( .A(n163), .Z(n186) );
  GTECH_XOR2 U164 ( .A(n187), .B(n165), .Z(n163) );
  GTECH_ADD_ABC U165 ( .A(n188), .B(n189), .C(n190), .COUT(n165) );
  GTECH_NOT U166 ( .A(n191), .Z(n190) );
  GTECH_XOR3 U167 ( .A(n192), .B(n193), .C(n194), .Z(n189) );
  GTECH_XNOR4 U168 ( .A(n170), .B(n183), .C(n168), .D(n169), .Z(n187) );
  GTECH_NOT U169 ( .A(n181), .Z(n169) );
  GTECH_OR_NOT U170 ( .A(n172), .B(I_a[6]), .Z(n181) );
  GTECH_XOR3 U171 ( .A(n176), .B(n178), .C(n177), .Z(n168) );
  GTECH_OAI21 U172 ( .A(n195), .B(n196), .C(n197), .Z(n177) );
  GTECH_OAI21 U173 ( .A(n198), .B(n199), .C(n200), .Z(n197) );
  GTECH_NOT U174 ( .A(n199), .Z(n195) );
  GTECH_NOT U175 ( .A(n201), .Z(n178) );
  GTECH_OR_NOT U176 ( .A(n202), .B(I_b[7]), .Z(n201) );
  GTECH_NOT U177 ( .A(n174), .Z(n176) );
  GTECH_OR_NOT U178 ( .A(n180), .B(I_b[6]), .Z(n174) );
  GTECH_OAI21 U179 ( .A(n194), .B(n203), .C(n204), .Z(n183) );
  GTECH_OAI21 U180 ( .A(n192), .B(n205), .C(n193), .Z(n204) );
  GTECH_NOT U181 ( .A(n205), .Z(n194) );
  GTECH_NOT U182 ( .A(n206), .Z(n170) );
  GTECH_OR_NOT U183 ( .A(n137), .B(I_a[5]), .Z(n206) );
  GTECH_NOT U184 ( .A(I_b[5]), .Z(n137) );
  GTECH_NOT U185 ( .A(n157), .Z(n161) );
  GTECH_XOR2 U186 ( .A(n185), .B(n154), .Z(n157) );
  GTECH_AOI2N2 U187 ( .A(n207), .B(n208), .C(n209), .D(n210), .Z(n154) );
  GTECH_OR_NOT U188 ( .A(n211), .B(n209), .Z(n208) );
  GTECH_XOR2 U189 ( .A(n212), .B(n153), .Z(n185) );
  GTECH_AND2 U190 ( .A(n213), .B(n214), .Z(n153) );
  GTECH_OR_NOT U191 ( .A(n215), .B(n216), .Z(n214) );
  GTECH_OAI21 U192 ( .A(n217), .B(n216), .C(n218), .Z(n213) );
  GTECH_OR_NOT U193 ( .A(n219), .B(I_a[7]), .Z(n212) );
  GTECH_NOT U194 ( .A(n162), .Z(n156) );
  GTECH_OAI2N2 U195 ( .A(n220), .B(n221), .C(n222), .D(n223), .Z(n162) );
  GTECH_OR_NOT U196 ( .A(n224), .B(n220), .Z(n223) );
  GTECH_XOR3 U197 ( .A(n220), .B(n224), .C(n225), .Z(N149) );
  GTECH_NOT U198 ( .A(n222), .Z(n225) );
  GTECH_XOR2 U199 ( .A(n226), .B(n188), .Z(n222) );
  GTECH_ADD_ABC U200 ( .A(n227), .B(n228), .C(n229), .COUT(n188) );
  GTECH_XOR3 U201 ( .A(n230), .B(n231), .C(n232), .Z(n228) );
  GTECH_OA21 U202 ( .A(n233), .B(n234), .C(n235), .Z(n227) );
  GTECH_XNOR4 U203 ( .A(n193), .B(n205), .C(n191), .D(n192), .Z(n226) );
  GTECH_NOT U204 ( .A(n203), .Z(n192) );
  GTECH_OR_NOT U205 ( .A(n172), .B(I_a[5]), .Z(n203) );
  GTECH_NOT U206 ( .A(I_b[4]), .Z(n172) );
  GTECH_XOR3 U207 ( .A(n198), .B(n200), .C(n199), .Z(n191) );
  GTECH_OAI21 U208 ( .A(n236), .B(n237), .C(n238), .Z(n199) );
  GTECH_NOT U209 ( .A(n239), .Z(n200) );
  GTECH_OR_NOT U210 ( .A(n240), .B(I_b[7]), .Z(n239) );
  GTECH_NOT U211 ( .A(n196), .Z(n198) );
  GTECH_OR_NOT U212 ( .A(n202), .B(I_b[6]), .Z(n196) );
  GTECH_OAI21 U213 ( .A(n232), .B(n241), .C(n242), .Z(n205) );
  GTECH_OAI21 U214 ( .A(n230), .B(n243), .C(n231), .Z(n242) );
  GTECH_NOT U215 ( .A(n243), .Z(n232) );
  GTECH_NOT U216 ( .A(n244), .Z(n193) );
  GTECH_OR_NOT U217 ( .A(n180), .B(I_b[5]), .Z(n244) );
  GTECH_NOT U218 ( .A(n221), .Z(n224) );
  GTECH_XOR3 U219 ( .A(n211), .B(n209), .C(n207), .Z(n221) );
  GTECH_XOR3 U220 ( .A(n217), .B(n218), .C(n216), .Z(n207) );
  GTECH_OAI21 U221 ( .A(n245), .B(n246), .C(n247), .Z(n216) );
  GTECH_OAI21 U222 ( .A(n248), .B(n249), .C(n250), .Z(n247) );
  GTECH_NOT U223 ( .A(n249), .Z(n245) );
  GTECH_NOT U224 ( .A(n251), .Z(n218) );
  GTECH_OR_NOT U225 ( .A(n219), .B(I_a[6]), .Z(n251) );
  GTECH_NOT U226 ( .A(n215), .Z(n217) );
  GTECH_OR_NOT U227 ( .A(n252), .B(I_a[7]), .Z(n215) );
  GTECH_ADD_ABC U228 ( .A(n253), .B(n254), .C(n255), .COUT(n209) );
  GTECH_XOR2 U229 ( .A(n256), .B(n257), .Z(n254) );
  GTECH_AND2 U230 ( .A(I_a[7]), .B(I_b[1]), .Z(n257) );
  GTECH_NOT U231 ( .A(n210), .Z(n211) );
  GTECH_OR_NOT U232 ( .A(n256), .B(I_a[7]), .Z(n210) );
  GTECH_ADD_ABC U233 ( .A(n258), .B(n259), .C(n260), .COUT(n220) );
  GTECH_XOR3 U234 ( .A(n253), .B(n261), .C(n255), .Z(n259) );
  GTECH_NOT U235 ( .A(n262), .Z(n255) );
  GTECH_XOR3 U236 ( .A(n263), .B(n260), .C(n258), .Z(N148) );
  GTECH_ADD_ABC U237 ( .A(n264), .B(n265), .C(n266), .COUT(n258) );
  GTECH_NOT U238 ( .A(n267), .Z(n266) );
  GTECH_XOR3 U239 ( .A(n268), .B(n269), .C(n270), .Z(n265) );
  GTECH_XOR2 U240 ( .A(n271), .B(n272), .Z(n260) );
  GTECH_OA21 U241 ( .A(n233), .B(n234), .C(n235), .Z(n272) );
  GTECH_OAI21 U242 ( .A(n273), .B(n274), .C(n275), .Z(n235) );
  GTECH_NOT U243 ( .A(n233), .Z(n274) );
  GTECH_XNOR4 U244 ( .A(n231), .B(n243), .C(n229), .D(n230), .Z(n271) );
  GTECH_NOT U245 ( .A(n241), .Z(n230) );
  GTECH_OR_NOT U246 ( .A(n180), .B(I_b[4]), .Z(n241) );
  GTECH_XOR3 U247 ( .A(n276), .B(n277), .C(n238), .Z(n229) );
  GTECH_NAND3 U248 ( .A(I_b[6]), .B(I_a[1]), .C(n278), .Z(n238) );
  GTECH_NOT U249 ( .A(n237), .Z(n277) );
  GTECH_OR_NOT U250 ( .A(n279), .B(I_b[7]), .Z(n237) );
  GTECH_NOT U251 ( .A(n236), .Z(n276) );
  GTECH_OR_NOT U252 ( .A(n240), .B(I_b[6]), .Z(n236) );
  GTECH_OAI21 U253 ( .A(n280), .B(n281), .C(n282), .Z(n243) );
  GTECH_OAI21 U254 ( .A(n283), .B(n284), .C(n285), .Z(n282) );
  GTECH_NOT U255 ( .A(n284), .Z(n280) );
  GTECH_NOT U256 ( .A(n286), .Z(n231) );
  GTECH_OR_NOT U257 ( .A(n202), .B(I_b[5]), .Z(n286) );
  GTECH_XOR3 U258 ( .A(n261), .B(n262), .C(n253), .Z(n263) );
  GTECH_ADD_ABC U259 ( .A(n268), .B(n287), .C(n270), .COUT(n253) );
  GTECH_NOT U260 ( .A(n288), .Z(n270) );
  GTECH_XOR3 U261 ( .A(n289), .B(n290), .C(n291), .Z(n287) );
  GTECH_XOR3 U262 ( .A(n248), .B(n250), .C(n249), .Z(n262) );
  GTECH_OAI21 U263 ( .A(n292), .B(n293), .C(n294), .Z(n249) );
  GTECH_OAI21 U264 ( .A(n295), .B(n296), .C(n297), .Z(n294) );
  GTECH_NOT U265 ( .A(n296), .Z(n292) );
  GTECH_NOT U266 ( .A(n298), .Z(n250) );
  GTECH_OR_NOT U267 ( .A(n219), .B(I_a[5]), .Z(n298) );
  GTECH_NOT U268 ( .A(I_b[3]), .Z(n219) );
  GTECH_NOT U269 ( .A(n246), .Z(n248) );
  GTECH_OR_NOT U270 ( .A(n252), .B(I_a[6]), .Z(n246) );
  GTECH_XOR2 U271 ( .A(n299), .B(n256), .Z(n261) );
  GTECH_OA21 U272 ( .A(n291), .B(n300), .C(n301), .Z(n256) );
  GTECH_OAI21 U273 ( .A(n289), .B(n302), .C(n290), .Z(n301) );
  GTECH_NOT U274 ( .A(n302), .Z(n291) );
  GTECH_AND2 U275 ( .A(I_b[1]), .B(I_a[7]), .Z(n299) );
  GTECH_XOR2 U276 ( .A(n303), .B(n264), .Z(N147) );
  GTECH_ADD_ABC U277 ( .A(n304), .B(n305), .C(n306), .COUT(n264) );
  GTECH_XOR3 U278 ( .A(n307), .B(n308), .C(n309), .Z(n305) );
  GTECH_NOT U279 ( .A(n310), .Z(n308) );
  GTECH_OA21 U280 ( .A(n311), .B(n312), .C(n313), .Z(n304) );
  GTECH_XNOR4 U281 ( .A(n269), .B(n288), .C(n267), .D(n268), .Z(n303) );
  GTECH_ADD_ABC U282 ( .A(n307), .B(n314), .C(n309), .COUT(n268) );
  GTECH_NOT U283 ( .A(n315), .Z(n309) );
  GTECH_XOR3 U284 ( .A(n316), .B(n317), .C(n318), .Z(n314) );
  GTECH_XOR3 U285 ( .A(n275), .B(n234), .C(n233), .Z(n267) );
  GTECH_XOR2 U286 ( .A(n319), .B(n278), .Z(n233) );
  GTECH_NOT U287 ( .A(n320), .Z(n278) );
  GTECH_OR_NOT U288 ( .A(n321), .B(I_b[7]), .Z(n320) );
  GTECH_OR_NOT U289 ( .A(n279), .B(I_b[6]), .Z(n319) );
  GTECH_NOT U290 ( .A(n273), .Z(n234) );
  GTECH_XOR3 U291 ( .A(n283), .B(n285), .C(n284), .Z(n273) );
  GTECH_OAI21 U292 ( .A(n322), .B(n323), .C(n324), .Z(n284) );
  GTECH_NOT U293 ( .A(n325), .Z(n285) );
  GTECH_OR_NOT U294 ( .A(n240), .B(I_b[5]), .Z(n325) );
  GTECH_NOT U295 ( .A(n281), .Z(n283) );
  GTECH_OR_NOT U296 ( .A(n202), .B(I_b[4]), .Z(n281) );
  GTECH_NOT U297 ( .A(n326), .Z(n275) );
  GTECH_NAND3 U298 ( .A(I_a[0]), .B(n327), .C(I_b[6]), .Z(n326) );
  GTECH_NOT U299 ( .A(n328), .Z(n327) );
  GTECH_XOR3 U300 ( .A(n295), .B(n297), .C(n296), .Z(n288) );
  GTECH_OAI21 U301 ( .A(n329), .B(n330), .C(n331), .Z(n296) );
  GTECH_OAI21 U302 ( .A(n332), .B(n333), .C(n334), .Z(n331) );
  GTECH_NOT U303 ( .A(n333), .Z(n329) );
  GTECH_NOT U304 ( .A(n335), .Z(n297) );
  GTECH_OR_NOT U305 ( .A(n180), .B(I_b[3]), .Z(n335) );
  GTECH_NOT U306 ( .A(n293), .Z(n295) );
  GTECH_OR_NOT U307 ( .A(n252), .B(I_a[5]), .Z(n293) );
  GTECH_NOT U308 ( .A(I_b[2]), .Z(n252) );
  GTECH_NOT U309 ( .A(n336), .Z(n269) );
  GTECH_XOR3 U310 ( .A(n289), .B(n290), .C(n302), .Z(n336) );
  GTECH_OAI21 U311 ( .A(n318), .B(n337), .C(n338), .Z(n302) );
  GTECH_OAI21 U312 ( .A(n316), .B(n339), .C(n317), .Z(n338) );
  GTECH_NOT U313 ( .A(n339), .Z(n318) );
  GTECH_NOT U314 ( .A(n340), .Z(n290) );
  GTECH_OR_NOT U315 ( .A(n341), .B(I_a[6]), .Z(n340) );
  GTECH_NOT U316 ( .A(n300), .Z(n289) );
  GTECH_OR_NOT U317 ( .A(n342), .B(I_a[7]), .Z(n300) );
  GTECH_XOR2 U318 ( .A(n343), .B(n344), .Z(N146) );
  GTECH_XNOR4 U319 ( .A(n315), .B(n307), .C(n310), .D(n306), .Z(n344) );
  GTECH_XOR2 U320 ( .A(n328), .B(n345), .Z(n306) );
  GTECH_AND2 U321 ( .A(I_b[6]), .B(I_a[0]), .Z(n345) );
  GTECH_XOR3 U322 ( .A(n346), .B(n347), .C(n324), .Z(n328) );
  GTECH_NAND3 U323 ( .A(I_b[4]), .B(I_a[1]), .C(n348), .Z(n324) );
  GTECH_NOT U324 ( .A(n323), .Z(n347) );
  GTECH_OR_NOT U325 ( .A(n279), .B(I_b[5]), .Z(n323) );
  GTECH_NOT U326 ( .A(n322), .Z(n346) );
  GTECH_OR_NOT U327 ( .A(n240), .B(I_b[4]), .Z(n322) );
  GTECH_XOR3 U328 ( .A(n316), .B(n317), .C(n339), .Z(n310) );
  GTECH_OAI21 U329 ( .A(n349), .B(n350), .C(n351), .Z(n339) );
  GTECH_OAI21 U330 ( .A(n352), .B(n353), .C(n354), .Z(n351) );
  GTECH_NOT U331 ( .A(n355), .Z(n317) );
  GTECH_OR_NOT U332 ( .A(n341), .B(I_a[5]), .Z(n355) );
  GTECH_NOT U333 ( .A(n337), .Z(n316) );
  GTECH_OR_NOT U334 ( .A(n342), .B(I_a[6]), .Z(n337) );
  GTECH_ADD_ABC U335 ( .A(n356), .B(n357), .C(n358), .COUT(n307) );
  GTECH_NOT U336 ( .A(n359), .Z(n358) );
  GTECH_XOR3 U337 ( .A(n352), .B(n354), .C(n349), .Z(n357) );
  GTECH_NOT U338 ( .A(n353), .Z(n349) );
  GTECH_XOR3 U339 ( .A(n332), .B(n334), .C(n333), .Z(n315) );
  GTECH_OAI21 U340 ( .A(n360), .B(n361), .C(n362), .Z(n333) );
  GTECH_OAI21 U341 ( .A(n363), .B(n364), .C(n365), .Z(n362) );
  GTECH_NOT U342 ( .A(n364), .Z(n360) );
  GTECH_NOT U343 ( .A(n366), .Z(n334) );
  GTECH_OR_NOT U344 ( .A(n202), .B(I_b[3]), .Z(n366) );
  GTECH_NOT U345 ( .A(n330), .Z(n332) );
  GTECH_OR_NOT U346 ( .A(n180), .B(I_b[2]), .Z(n330) );
  GTECH_NOT U347 ( .A(I_a[4]), .Z(n180) );
  GTECH_OA21 U348 ( .A(n311), .B(n312), .C(n313), .Z(n343) );
  GTECH_OAI21 U349 ( .A(n367), .B(n368), .C(n369), .Z(n313) );
  GTECH_NOT U350 ( .A(n311), .Z(n368) );
  GTECH_XOR3 U351 ( .A(n369), .B(n312), .C(n311), .Z(N145) );
  GTECH_XOR2 U352 ( .A(n370), .B(n348), .Z(n311) );
  GTECH_NOT U353 ( .A(n371), .Z(n348) );
  GTECH_OR_NOT U354 ( .A(n321), .B(I_b[5]), .Z(n371) );
  GTECH_OR_NOT U355 ( .A(n279), .B(I_b[4]), .Z(n370) );
  GTECH_NOT U356 ( .A(n367), .Z(n312) );
  GTECH_XOR2 U357 ( .A(n372), .B(n356), .Z(n367) );
  GTECH_ADD_ABC U358 ( .A(n373), .B(n374), .C(n375), .COUT(n356) );
  GTECH_XOR3 U359 ( .A(n376), .B(n377), .C(n378), .Z(n374) );
  GTECH_OA21 U360 ( .A(n379), .B(n380), .C(n381), .Z(n373) );
  GTECH_XNOR4 U361 ( .A(n354), .B(n353), .C(n359), .D(n352), .Z(n372) );
  GTECH_NOT U362 ( .A(n350), .Z(n352) );
  GTECH_OR_NOT U363 ( .A(n342), .B(I_a[5]), .Z(n350) );
  GTECH_XOR3 U364 ( .A(n363), .B(n365), .C(n364), .Z(n359) );
  GTECH_OAI21 U365 ( .A(n382), .B(n383), .C(n384), .Z(n364) );
  GTECH_NOT U366 ( .A(n385), .Z(n365) );
  GTECH_OR_NOT U367 ( .A(n240), .B(I_b[3]), .Z(n385) );
  GTECH_NOT U368 ( .A(n361), .Z(n363) );
  GTECH_OR_NOT U369 ( .A(n202), .B(I_b[2]), .Z(n361) );
  GTECH_OAI21 U370 ( .A(n378), .B(n386), .C(n387), .Z(n353) );
  GTECH_OAI21 U371 ( .A(n376), .B(n388), .C(n377), .Z(n387) );
  GTECH_NOT U372 ( .A(n386), .Z(n376) );
  GTECH_NOT U373 ( .A(n388), .Z(n378) );
  GTECH_NOT U374 ( .A(n389), .Z(n354) );
  GTECH_OR_NOT U375 ( .A(n341), .B(I_a[4]), .Z(n389) );
  GTECH_NOT U376 ( .A(n390), .Z(n369) );
  GTECH_NAND3 U377 ( .A(I_a[0]), .B(n391), .C(I_b[4]), .Z(n390) );
  GTECH_XOR2 U378 ( .A(n392), .B(n391), .Z(N144) );
  GTECH_XOR2 U379 ( .A(n393), .B(n394), .Z(n391) );
  GTECH_XNOR4 U380 ( .A(n377), .B(n388), .C(n386), .D(n375), .Z(n394) );
  GTECH_XOR3 U381 ( .A(n395), .B(n396), .C(n384), .Z(n375) );
  GTECH_NAND3 U382 ( .A(I_b[2]), .B(I_a[1]), .C(n397), .Z(n384) );
  GTECH_NOT U383 ( .A(n383), .Z(n396) );
  GTECH_OR_NOT U384 ( .A(n279), .B(I_b[3]), .Z(n383) );
  GTECH_NOT U385 ( .A(n382), .Z(n395) );
  GTECH_OR_NOT U386 ( .A(n240), .B(I_b[2]), .Z(n382) );
  GTECH_OR_NOT U387 ( .A(n342), .B(I_a[4]), .Z(n386) );
  GTECH_NOT U388 ( .A(I_b[0]), .Z(n342) );
  GTECH_OAI21 U389 ( .A(n398), .B(n399), .C(n400), .Z(n388) );
  GTECH_OAI21 U390 ( .A(n401), .B(n402), .C(n403), .Z(n400) );
  GTECH_NOT U391 ( .A(n402), .Z(n398) );
  GTECH_NOT U392 ( .A(n404), .Z(n377) );
  GTECH_OR_NOT U393 ( .A(n341), .B(I_a[3]), .Z(n404) );
  GTECH_OA21 U394 ( .A(n379), .B(n380), .C(n381), .Z(n393) );
  GTECH_OAI21 U395 ( .A(n405), .B(n406), .C(n407), .Z(n381) );
  GTECH_NOT U396 ( .A(n379), .Z(n406) );
  GTECH_AND2 U397 ( .A(I_b[4]), .B(I_a[0]), .Z(n392) );
  GTECH_XOR3 U398 ( .A(n407), .B(n380), .C(n379), .Z(N143) );
  GTECH_XOR2 U399 ( .A(n408), .B(n397), .Z(n379) );
  GTECH_NOT U400 ( .A(n409), .Z(n397) );
  GTECH_OR_NOT U401 ( .A(n321), .B(I_b[3]), .Z(n409) );
  GTECH_NOT U402 ( .A(I_a[0]), .Z(n321) );
  GTECH_OR_NOT U403 ( .A(n279), .B(I_b[2]), .Z(n408) );
  GTECH_NOT U404 ( .A(I_a[1]), .Z(n279) );
  GTECH_NOT U405 ( .A(n405), .Z(n380) );
  GTECH_XOR3 U406 ( .A(n401), .B(n403), .C(n402), .Z(n405) );
  GTECH_OAI21 U407 ( .A(n410), .B(n411), .C(n412), .Z(n402) );
  GTECH_NOT U408 ( .A(n413), .Z(n403) );
  GTECH_OR_NOT U409 ( .A(n240), .B(I_b[1]), .Z(n413) );
  GTECH_NOT U410 ( .A(n399), .Z(n401) );
  GTECH_OR_NOT U411 ( .A(n202), .B(I_b[0]), .Z(n399) );
  GTECH_NOT U412 ( .A(I_a[3]), .Z(n202) );
  GTECH_NOT U413 ( .A(n414), .Z(n407) );
  GTECH_NAND3 U414 ( .A(I_a[0]), .B(n415), .C(I_b[2]), .Z(n414) );
  GTECH_XOR2 U415 ( .A(n416), .B(n415), .Z(N142) );
  GTECH_NOT U416 ( .A(n417), .Z(n415) );
  GTECH_XOR3 U417 ( .A(n418), .B(n419), .C(n412), .Z(n417) );
  GTECH_NAND3 U418 ( .A(n420), .B(I_b[0]), .C(I_a[1]), .Z(n412) );
  GTECH_NOT U419 ( .A(n410), .Z(n419) );
  GTECH_OR_NOT U420 ( .A(n341), .B(I_a[1]), .Z(n410) );
  GTECH_NOT U421 ( .A(n411), .Z(n418) );
  GTECH_OR_NOT U422 ( .A(n240), .B(I_b[0]), .Z(n411) );
  GTECH_NOT U423 ( .A(I_a[2]), .Z(n240) );
  GTECH_AND2 U424 ( .A(I_b[2]), .B(I_a[0]), .Z(n416) );
  GTECH_XOR2 U425 ( .A(n420), .B(n421), .Z(N141) );
  GTECH_AND2 U426 ( .A(I_a[1]), .B(I_b[0]), .Z(n421) );
  GTECH_NOT U427 ( .A(n422), .Z(n420) );
  GTECH_OR_NOT U428 ( .A(n341), .B(I_a[0]), .Z(n422) );
  GTECH_NOT U429 ( .A(I_b[1]), .Z(n341) );
  GTECH_AND2 U430 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

