
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121;

  GTECH_XOR2 U81 ( .A(n62), .B(n63), .Z(sum[9]) );
  GTECH_XOR2 U82 ( .A(n64), .B(n65), .Z(sum[8]) );
  GTECH_XNOR2 U83 ( .A(n66), .B(n67), .Z(sum[7]) );
  GTECH_AOI21 U84 ( .A(n68), .B(n69), .C(n70), .Z(n67) );
  GTECH_XOR2 U85 ( .A(n69), .B(n68), .Z(sum[6]) );
  GTECH_AO22 U86 ( .A(b[5]), .B(a[5]), .C(n71), .D(n72), .Z(n68) );
  GTECH_XOR2 U87 ( .A(n72), .B(n71), .Z(sum[5]) );
  GTECH_AO22 U88 ( .A(n73), .B(n74), .C(b[4]), .D(a[4]), .Z(n71) );
  GTECH_XOR2 U89 ( .A(n74), .B(n73), .Z(sum[4]) );
  GTECH_XNOR2 U90 ( .A(n75), .B(n76), .Z(sum[3]) );
  GTECH_AOI21 U91 ( .A(n77), .B(n78), .C(n79), .Z(n76) );
  GTECH_XOR2 U92 ( .A(n77), .B(n78), .Z(sum[2]) );
  GTECH_AO21 U93 ( .A(n80), .B(n81), .C(n82), .Z(n77) );
  GTECH_XOR2 U94 ( .A(n81), .B(n80), .Z(sum[1]) );
  GTECH_AO21 U95 ( .A(cin), .B(n83), .C(n84), .Z(n81) );
  GTECH_XNOR2 U96 ( .A(n85), .B(n86), .Z(sum[15]) );
  GTECH_AOI21 U97 ( .A(n87), .B(n88), .C(n89), .Z(n86) );
  GTECH_XOR2 U98 ( .A(n88), .B(n87), .Z(sum[14]) );
  GTECH_AO22 U99 ( .A(n90), .B(n91), .C(b[13]), .D(a[13]), .Z(n87) );
  GTECH_XOR2 U100 ( .A(n91), .B(n90), .Z(sum[13]) );
  GTECH_AO22 U101 ( .A(a[12]), .B(b[12]), .C(cout), .D(n92), .Z(n90) );
  GTECH_XOR2 U102 ( .A(n92), .B(cout), .Z(sum[12]) );
  GTECH_XNOR2 U103 ( .A(n93), .B(n94), .Z(sum[11]) );
  GTECH_AOI21 U104 ( .A(n95), .B(n96), .C(n97), .Z(n94) );
  GTECH_XOR2 U105 ( .A(n96), .B(n95), .Z(sum[10]) );
  GTECH_AO22 U106 ( .A(n63), .B(n62), .C(b[9]), .D(a[9]), .Z(n95) );
  GTECH_AO22 U107 ( .A(a[8]), .B(b[8]), .C(n65), .D(n64), .Z(n63) );
  GTECH_XOR2 U108 ( .A(cin), .B(n83), .Z(sum[0]) );
  GTECH_AO21 U109 ( .A(n98), .B(n65), .C(n99), .Z(cout) );
  GTECH_AO21 U110 ( .A(n100), .B(n73), .C(n101), .Z(n65) );
  GTECH_AO21 U111 ( .A(cin), .B(n102), .C(n103), .Z(n73) );
  GTECH_AND3 U112 ( .A(n100), .B(n102), .C(n98), .Z(Pm) );
  GTECH_AND5 U113 ( .A(n80), .B(n75), .C(n78), .D(n83), .E(n104), .Z(n102) );
  GTECH_OA21 U114 ( .A(b[0]), .B(a[0]), .C(n105), .Z(n83) );
  GTECH_NOT U115 ( .A(n84), .Z(n105) );
  GTECH_AO21 U116 ( .A(n98), .B(n106), .C(n99), .Z(Gm) );
  GTECH_AO22 U117 ( .A(b[15]), .B(a[15]), .C(n107), .D(n85), .Z(n99) );
  GTECH_AO21 U118 ( .A(n108), .B(n88), .C(n89), .Z(n107) );
  GTECH_AND2 U119 ( .A(a[14]), .B(b[14]), .Z(n89) );
  GTECH_AO21 U120 ( .A(b[13]), .B(a[13]), .C(n109), .Z(n108) );
  GTECH_AND3 U121 ( .A(a[12]), .B(n91), .C(b[12]), .Z(n109) );
  GTECH_AO21 U122 ( .A(n100), .B(n103), .C(n101), .Z(n106) );
  GTECH_AO22 U123 ( .A(b[11]), .B(a[11]), .C(n110), .D(n93), .Z(n101) );
  GTECH_AO21 U124 ( .A(n111), .B(n96), .C(n97), .Z(n110) );
  GTECH_AND2 U125 ( .A(a[10]), .B(b[10]), .Z(n97) );
  GTECH_AO21 U126 ( .A(b[9]), .B(a[9]), .C(n112), .Z(n111) );
  GTECH_AND3 U127 ( .A(a[8]), .B(n62), .C(b[8]), .Z(n112) );
  GTECH_NOT U128 ( .A(n113), .Z(n103) );
  GTECH_AOI222 U129 ( .A(a[7]), .B(b[7]), .C(n104), .D(n114), .E(n66), .F(n115), .Z(n113) );
  GTECH_AO21 U130 ( .A(n69), .B(n116), .C(n70), .Z(n115) );
  GTECH_AND2 U131 ( .A(a[6]), .B(b[6]), .Z(n70) );
  GTECH_AO22 U132 ( .A(a[4]), .B(n117), .C(b[5]), .D(a[5]), .Z(n116) );
  GTECH_AND2 U133 ( .A(n72), .B(b[4]), .Z(n117) );
  GTECH_AO22 U134 ( .A(n118), .B(n75), .C(b[3]), .D(a[3]), .Z(n114) );
  GTECH_XOR2 U135 ( .A(a[3]), .B(b[3]), .Z(n75) );
  GTECH_AO21 U136 ( .A(n119), .B(n78), .C(n79), .Z(n118) );
  GTECH_OA21 U137 ( .A(b[2]), .B(a[2]), .C(n120), .Z(n78) );
  GTECH_NOT U138 ( .A(n79), .Z(n120) );
  GTECH_AND2 U139 ( .A(a[2]), .B(b[2]), .Z(n79) );
  GTECH_AO21 U140 ( .A(n84), .B(n80), .C(n82), .Z(n119) );
  GTECH_OA21 U141 ( .A(b[1]), .B(a[1]), .C(n121), .Z(n80) );
  GTECH_NOT U142 ( .A(n82), .Z(n121) );
  GTECH_AND2 U143 ( .A(a[1]), .B(b[1]), .Z(n82) );
  GTECH_AND2 U144 ( .A(b[0]), .B(a[0]), .Z(n84) );
  GTECH_AND4 U145 ( .A(n74), .B(n72), .C(n69), .D(n66), .Z(n104) );
  GTECH_XOR2 U146 ( .A(a[7]), .B(b[7]), .Z(n66) );
  GTECH_XOR2 U147 ( .A(a[6]), .B(b[6]), .Z(n69) );
  GTECH_XOR2 U148 ( .A(a[5]), .B(b[5]), .Z(n72) );
  GTECH_XOR2 U149 ( .A(a[4]), .B(b[4]), .Z(n74) );
  GTECH_AND4 U150 ( .A(n64), .B(n93), .C(n96), .D(n62), .Z(n100) );
  GTECH_XOR2 U151 ( .A(a[9]), .B(b[9]), .Z(n62) );
  GTECH_XOR2 U152 ( .A(a[10]), .B(b[10]), .Z(n96) );
  GTECH_XOR2 U153 ( .A(a[11]), .B(b[11]), .Z(n93) );
  GTECH_XOR2 U154 ( .A(a[8]), .B(b[8]), .Z(n64) );
  GTECH_AND4 U155 ( .A(n92), .B(n85), .C(n88), .D(n91), .Z(n98) );
  GTECH_XOR2 U156 ( .A(a[13]), .B(b[13]), .Z(n91) );
  GTECH_XOR2 U157 ( .A(a[14]), .B(b[14]), .Z(n88) );
  GTECH_XOR2 U158 ( .A(a[15]), .B(b[15]), .Z(n85) );
  GTECH_XOR2 U159 ( .A(a[12]), .B(b[12]), .Z(n92) );
endmodule

