
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_OAI21 U75 ( .A(n83), .B(n84), .C(n85), .Z(N155) );
  GTECH_OA22 U76 ( .A(n86), .B(n87), .C(n88), .D(n89), .Z(n85) );
  GTECH_NOT U77 ( .A(n90), .Z(n87) );
  GTECH_XOR2 U78 ( .A(n91), .B(n92), .Z(N154) );
  GTECH_NOT U79 ( .A(n83), .Z(n92) );
  GTECH_XOR2 U80 ( .A(n90), .B(n86), .Z(n83) );
  GTECH_AOI2N2 U81 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n86) );
  GTECH_NAND2 U82 ( .A(n95), .B(n96), .Z(n94) );
  GTECH_XOR2 U83 ( .A(n89), .B(n88), .Z(n90) );
  GTECH_OA21 U84 ( .A(n97), .B(n98), .C(n99), .Z(n88) );
  GTECH_OAI21 U85 ( .A(n100), .B(n101), .C(n102), .Z(n99) );
  GTECH_NAND2 U86 ( .A(I_b[7]), .B(I_a[7]), .Z(n89) );
  GTECH_NOT U87 ( .A(n84), .Z(n91) );
  GTECH_NAND2 U88 ( .A(n103), .B(n104), .Z(n84) );
  GTECH_XOR2 U89 ( .A(n104), .B(n103), .Z(N153) );
  GTECH_NOT U90 ( .A(n105), .Z(n103) );
  GTECH_XNOR3 U91 ( .A(n106), .B(n95), .C(n107), .Z(n105) );
  GTECH_NOT U92 ( .A(n93), .Z(n107) );
  GTECH_XNOR3 U93 ( .A(n100), .B(n102), .C(n97), .Z(n93) );
  GTECH_NOT U94 ( .A(n101), .Z(n97) );
  GTECH_OAI21 U95 ( .A(n108), .B(n109), .C(n110), .Z(n101) );
  GTECH_OAI21 U96 ( .A(n111), .B(n112), .C(n113), .Z(n110) );
  GTECH_NOT U97 ( .A(n114), .Z(n102) );
  GTECH_NAND2 U98 ( .A(I_b[7]), .B(I_a[6]), .Z(n114) );
  GTECH_NOT U99 ( .A(n98), .Z(n100) );
  GTECH_NAND2 U100 ( .A(I_a[7]), .B(I_b[6]), .Z(n98) );
  GTECH_ADD_ABC U101 ( .A(n115), .B(n116), .C(n117), .COUT(n95) );
  GTECH_NOT U102 ( .A(n118), .Z(n117) );
  GTECH_XOR2 U103 ( .A(n119), .B(n120), .Z(n116) );
  GTECH_AND2 U104 ( .A(I_a[7]), .B(I_b[5]), .Z(n120) );
  GTECH_NOT U105 ( .A(n96), .Z(n106) );
  GTECH_NAND2 U106 ( .A(I_a[7]), .B(n121), .Z(n96) );
  GTECH_NOT U107 ( .A(n122), .Z(n104) );
  GTECH_NAND2 U108 ( .A(n123), .B(n124), .Z(n122) );
  GTECH_NOT U109 ( .A(n125), .Z(n124) );
  GTECH_XOR2 U110 ( .A(n125), .B(n126), .Z(N152) );
  GTECH_NOT U111 ( .A(n123), .Z(n126) );
  GTECH_XOR4 U112 ( .A(n127), .B(n119), .C(n118), .D(n115), .Z(n123) );
  GTECH_ADD_ABC U113 ( .A(n128), .B(n129), .C(n130), .COUT(n115) );
  GTECH_XNOR3 U114 ( .A(n131), .B(n132), .C(n133), .Z(n129) );
  GTECH_XNOR3 U115 ( .A(n111), .B(n113), .C(n108), .Z(n118) );
  GTECH_NOT U116 ( .A(n112), .Z(n108) );
  GTECH_OAI21 U117 ( .A(n134), .B(n135), .C(n136), .Z(n112) );
  GTECH_OAI21 U118 ( .A(n137), .B(n138), .C(n139), .Z(n136) );
  GTECH_NOT U119 ( .A(n140), .Z(n113) );
  GTECH_NAND2 U120 ( .A(I_b[7]), .B(I_a[5]), .Z(n140) );
  GTECH_NOT U121 ( .A(n109), .Z(n111) );
  GTECH_NAND2 U122 ( .A(I_b[6]), .B(I_a[6]), .Z(n109) );
  GTECH_NOT U123 ( .A(n121), .Z(n119) );
  GTECH_OAI21 U124 ( .A(n141), .B(n142), .C(n143), .Z(n121) );
  GTECH_OAI21 U125 ( .A(n131), .B(n133), .C(n132), .Z(n143) );
  GTECH_AND2 U126 ( .A(I_a[7]), .B(I_b[5]), .Z(n127) );
  GTECH_ADD_ABC U127 ( .A(n144), .B(n145), .C(n146), .COUT(n125) );
  GTECH_OA22 U128 ( .A(n147), .B(n148), .C(n149), .D(n150), .Z(n145) );
  GTECH_OA21 U129 ( .A(n151), .B(n152), .C(n153), .Z(n144) );
  GTECH_XNOR3 U130 ( .A(n154), .B(n146), .C(n155), .Z(N151) );
  GTECH_OA21 U131 ( .A(n151), .B(n152), .C(n153), .Z(n155) );
  GTECH_OAI21 U132 ( .A(n156), .B(n157), .C(n158), .Z(n153) );
  GTECH_XOR2 U133 ( .A(n128), .B(n159), .Z(n146) );
  GTECH_XOR4 U134 ( .A(n132), .B(n141), .C(n130), .D(n131), .Z(n159) );
  GTECH_NOT U135 ( .A(n142), .Z(n131) );
  GTECH_NAND2 U136 ( .A(I_a[7]), .B(I_b[4]), .Z(n142) );
  GTECH_NOT U137 ( .A(n160), .Z(n130) );
  GTECH_XNOR3 U138 ( .A(n137), .B(n139), .C(n134), .Z(n160) );
  GTECH_NOT U139 ( .A(n138), .Z(n134) );
  GTECH_OAI21 U140 ( .A(n161), .B(n162), .C(n163), .Z(n138) );
  GTECH_OAI21 U141 ( .A(n164), .B(n165), .C(n166), .Z(n163) );
  GTECH_NOT U142 ( .A(n167), .Z(n139) );
  GTECH_NAND2 U143 ( .A(I_b[7]), .B(I_a[4]), .Z(n167) );
  GTECH_NOT U144 ( .A(n135), .Z(n137) );
  GTECH_NAND2 U145 ( .A(I_b[6]), .B(I_a[5]), .Z(n135) );
  GTECH_NOT U146 ( .A(n133), .Z(n141) );
  GTECH_OAI21 U147 ( .A(n168), .B(n169), .C(n170), .Z(n133) );
  GTECH_OAI21 U148 ( .A(n171), .B(n172), .C(n173), .Z(n170) );
  GTECH_NOT U149 ( .A(n174), .Z(n132) );
  GTECH_NAND2 U150 ( .A(I_a[6]), .B(I_b[5]), .Z(n174) );
  GTECH_ADD_ABC U151 ( .A(n175), .B(n176), .C(n177), .COUT(n128) );
  GTECH_NOT U152 ( .A(n178), .Z(n177) );
  GTECH_XNOR3 U153 ( .A(n171), .B(n173), .C(n172), .Z(n176) );
  GTECH_OA22 U154 ( .A(n147), .B(n148), .C(n149), .D(n150), .Z(n154) );
  GTECH_NOT U155 ( .A(n179), .Z(n150) );
  GTECH_NOT U156 ( .A(I_a[7]), .Z(n148) );
  GTECH_XNOR3 U157 ( .A(n151), .B(n156), .C(n158), .Z(N150) );
  GTECH_XOR2 U158 ( .A(n180), .B(n175), .Z(n158) );
  GTECH_ADD_ABC U159 ( .A(n181), .B(n182), .C(n183), .COUT(n175) );
  GTECH_NOT U160 ( .A(n184), .Z(n183) );
  GTECH_XNOR3 U161 ( .A(n185), .B(n186), .C(n187), .Z(n182) );
  GTECH_XOR4 U162 ( .A(n173), .B(n168), .C(n178), .D(n171), .Z(n180) );
  GTECH_NOT U163 ( .A(n169), .Z(n171) );
  GTECH_NAND2 U164 ( .A(I_a[6]), .B(I_b[4]), .Z(n169) );
  GTECH_XNOR3 U165 ( .A(n164), .B(n166), .C(n161), .Z(n178) );
  GTECH_NOT U166 ( .A(n165), .Z(n161) );
  GTECH_OAI21 U167 ( .A(n188), .B(n189), .C(n190), .Z(n165) );
  GTECH_OAI21 U168 ( .A(n191), .B(n192), .C(n193), .Z(n190) );
  GTECH_NOT U169 ( .A(n194), .Z(n166) );
  GTECH_NAND2 U170 ( .A(I_b[7]), .B(I_a[3]), .Z(n194) );
  GTECH_NOT U171 ( .A(n162), .Z(n164) );
  GTECH_NAND2 U172 ( .A(I_b[6]), .B(I_a[4]), .Z(n162) );
  GTECH_NOT U173 ( .A(n172), .Z(n168) );
  GTECH_OAI21 U174 ( .A(n195), .B(n196), .C(n197), .Z(n172) );
  GTECH_OAI21 U175 ( .A(n185), .B(n187), .C(n186), .Z(n197) );
  GTECH_NOT U176 ( .A(n198), .Z(n173) );
  GTECH_NAND2 U177 ( .A(I_a[5]), .B(I_b[5]), .Z(n198) );
  GTECH_NOT U178 ( .A(n152), .Z(n156) );
  GTECH_XOR2 U179 ( .A(n179), .B(n149), .Z(n152) );
  GTECH_AOI2N2 U180 ( .A(n199), .B(n200), .C(n201), .D(n202), .Z(n149) );
  GTECH_NAND2 U181 ( .A(n201), .B(n202), .Z(n200) );
  GTECH_XOR2 U182 ( .A(n203), .B(n147), .Z(n179) );
  GTECH_OA21 U183 ( .A(n204), .B(n205), .C(n206), .Z(n147) );
  GTECH_OAI21 U184 ( .A(n207), .B(n208), .C(n209), .Z(n206) );
  GTECH_NAND2 U185 ( .A(I_a[7]), .B(I_b[3]), .Z(n203) );
  GTECH_NOT U186 ( .A(n157), .Z(n151) );
  GTECH_OAI2N2 U187 ( .A(n210), .B(n211), .C(n212), .D(n213), .Z(n157) );
  GTECH_NAND2 U188 ( .A(n210), .B(n211), .Z(n213) );
  GTECH_XNOR3 U189 ( .A(n210), .B(n214), .C(n212), .Z(N149) );
  GTECH_XOR2 U190 ( .A(n215), .B(n181), .Z(n212) );
  GTECH_ADD_ABC U191 ( .A(n216), .B(n217), .C(n218), .COUT(n181) );
  GTECH_XNOR3 U192 ( .A(n219), .B(n220), .C(n221), .Z(n217) );
  GTECH_OA21 U193 ( .A(n222), .B(n223), .C(n224), .Z(n216) );
  GTECH_XOR4 U194 ( .A(n186), .B(n195), .C(n184), .D(n185), .Z(n215) );
  GTECH_NOT U195 ( .A(n196), .Z(n185) );
  GTECH_NAND2 U196 ( .A(I_a[5]), .B(I_b[4]), .Z(n196) );
  GTECH_XNOR3 U197 ( .A(n191), .B(n193), .C(n188), .Z(n184) );
  GTECH_NOT U198 ( .A(n192), .Z(n188) );
  GTECH_OAI21 U199 ( .A(n225), .B(n226), .C(n227), .Z(n192) );
  GTECH_NOT U200 ( .A(n228), .Z(n193) );
  GTECH_NAND2 U201 ( .A(I_b[7]), .B(I_a[2]), .Z(n228) );
  GTECH_NOT U202 ( .A(n189), .Z(n191) );
  GTECH_NAND2 U203 ( .A(I_b[6]), .B(I_a[3]), .Z(n189) );
  GTECH_NOT U204 ( .A(n187), .Z(n195) );
  GTECH_OAI21 U205 ( .A(n229), .B(n230), .C(n231), .Z(n187) );
  GTECH_OAI21 U206 ( .A(n219), .B(n221), .C(n220), .Z(n231) );
  GTECH_NOT U207 ( .A(n232), .Z(n186) );
  GTECH_NAND2 U208 ( .A(I_b[5]), .B(I_a[4]), .Z(n232) );
  GTECH_NOT U209 ( .A(n211), .Z(n214) );
  GTECH_XNOR3 U210 ( .A(n233), .B(n201), .C(n234), .Z(n211) );
  GTECH_NOT U211 ( .A(n199), .Z(n234) );
  GTECH_XNOR3 U212 ( .A(n207), .B(n209), .C(n204), .Z(n199) );
  GTECH_NOT U213 ( .A(n208), .Z(n204) );
  GTECH_OAI21 U214 ( .A(n235), .B(n236), .C(n237), .Z(n208) );
  GTECH_OAI21 U215 ( .A(n238), .B(n239), .C(n240), .Z(n237) );
  GTECH_NOT U216 ( .A(n241), .Z(n209) );
  GTECH_NAND2 U217 ( .A(I_a[6]), .B(I_b[3]), .Z(n241) );
  GTECH_NOT U218 ( .A(n205), .Z(n207) );
  GTECH_NAND2 U219 ( .A(I_a[7]), .B(I_b[2]), .Z(n205) );
  GTECH_ADD_ABC U220 ( .A(n242), .B(n243), .C(n244), .COUT(n201) );
  GTECH_NOT U221 ( .A(n245), .Z(n244) );
  GTECH_XOR2 U222 ( .A(n246), .B(n247), .Z(n243) );
  GTECH_AND2 U223 ( .A(I_a[7]), .B(I_b[1]), .Z(n247) );
  GTECH_NOT U224 ( .A(n202), .Z(n233) );
  GTECH_NAND2 U225 ( .A(I_a[7]), .B(n248), .Z(n202) );
  GTECH_ADD_ABC U226 ( .A(n249), .B(n250), .C(n251), .COUT(n210) );
  GTECH_XNOR3 U227 ( .A(n242), .B(n252), .C(n245), .Z(n250) );
  GTECH_XOR2 U228 ( .A(n253), .B(n249), .Z(N148) );
  GTECH_ADD_ABC U229 ( .A(n254), .B(n255), .C(n256), .COUT(n249) );
  GTECH_NOT U230 ( .A(n257), .Z(n256) );
  GTECH_XNOR3 U231 ( .A(n258), .B(n259), .C(n260), .Z(n255) );
  GTECH_XOR4 U232 ( .A(n252), .B(n242), .C(n245), .D(n251), .Z(n253) );
  GTECH_XOR2 U233 ( .A(n261), .B(n262), .Z(n251) );
  GTECH_XOR4 U234 ( .A(n220), .B(n229), .C(n218), .D(n219), .Z(n262) );
  GTECH_NOT U235 ( .A(n230), .Z(n219) );
  GTECH_NAND2 U236 ( .A(I_b[4]), .B(I_a[4]), .Z(n230) );
  GTECH_XNOR3 U237 ( .A(n263), .B(n264), .C(n265), .Z(n218) );
  GTECH_NOT U238 ( .A(n227), .Z(n265) );
  GTECH_NAND3 U239 ( .A(I_b[6]), .B(I_a[1]), .C(n266), .Z(n227) );
  GTECH_NOT U240 ( .A(n226), .Z(n264) );
  GTECH_NAND2 U241 ( .A(I_b[7]), .B(I_a[1]), .Z(n226) );
  GTECH_NOT U242 ( .A(n225), .Z(n263) );
  GTECH_NAND2 U243 ( .A(I_b[6]), .B(I_a[2]), .Z(n225) );
  GTECH_NOT U244 ( .A(n221), .Z(n229) );
  GTECH_OAI21 U245 ( .A(n267), .B(n268), .C(n269), .Z(n221) );
  GTECH_OAI21 U246 ( .A(n270), .B(n271), .C(n272), .Z(n269) );
  GTECH_NOT U247 ( .A(n273), .Z(n220) );
  GTECH_NAND2 U248 ( .A(I_b[5]), .B(I_a[3]), .Z(n273) );
  GTECH_OA21 U249 ( .A(n222), .B(n223), .C(n224), .Z(n261) );
  GTECH_OAI21 U250 ( .A(n274), .B(n275), .C(n276), .Z(n224) );
  GTECH_XNOR3 U251 ( .A(n238), .B(n240), .C(n235), .Z(n245) );
  GTECH_NOT U252 ( .A(n239), .Z(n235) );
  GTECH_OAI21 U253 ( .A(n277), .B(n278), .C(n279), .Z(n239) );
  GTECH_OAI21 U254 ( .A(n280), .B(n281), .C(n282), .Z(n279) );
  GTECH_NOT U255 ( .A(n283), .Z(n240) );
  GTECH_NAND2 U256 ( .A(I_a[5]), .B(I_b[3]), .Z(n283) );
  GTECH_NOT U257 ( .A(n236), .Z(n238) );
  GTECH_NAND2 U258 ( .A(I_a[6]), .B(I_b[2]), .Z(n236) );
  GTECH_ADD_ABC U259 ( .A(n258), .B(n284), .C(n285), .COUT(n242) );
  GTECH_XNOR3 U260 ( .A(n286), .B(n287), .C(n288), .Z(n284) );
  GTECH_XOR2 U261 ( .A(n289), .B(n246), .Z(n252) );
  GTECH_NOT U262 ( .A(n248), .Z(n246) );
  GTECH_OAI21 U263 ( .A(n290), .B(n291), .C(n292), .Z(n248) );
  GTECH_OAI21 U264 ( .A(n286), .B(n288), .C(n287), .Z(n292) );
  GTECH_AND2 U265 ( .A(I_a[7]), .B(I_b[1]), .Z(n289) );
  GTECH_XOR2 U266 ( .A(n293), .B(n254), .Z(N147) );
  GTECH_ADD_ABC U267 ( .A(n294), .B(n295), .C(n296), .COUT(n254) );
  GTECH_XNOR3 U268 ( .A(n297), .B(n298), .C(n299), .Z(n295) );
  GTECH_OA21 U269 ( .A(n300), .B(n301), .C(n302), .Z(n294) );
  GTECH_XOR4 U270 ( .A(n259), .B(n285), .C(n257), .D(n258), .Z(n293) );
  GTECH_ADD_ABC U271 ( .A(n297), .B(n303), .C(n304), .COUT(n258) );
  GTECH_NOT U272 ( .A(n299), .Z(n304) );
  GTECH_XNOR3 U273 ( .A(n305), .B(n306), .C(n307), .Z(n303) );
  GTECH_XNOR3 U274 ( .A(n276), .B(n223), .C(n275), .Z(n257) );
  GTECH_NOT U275 ( .A(n222), .Z(n275) );
  GTECH_XOR2 U276 ( .A(n308), .B(n266), .Z(n222) );
  GTECH_NOT U277 ( .A(n309), .Z(n266) );
  GTECH_NAND2 U278 ( .A(I_b[7]), .B(I_a[0]), .Z(n309) );
  GTECH_NAND2 U279 ( .A(I_b[6]), .B(I_a[1]), .Z(n308) );
  GTECH_NOT U280 ( .A(n274), .Z(n223) );
  GTECH_XNOR3 U281 ( .A(n270), .B(n272), .C(n267), .Z(n274) );
  GTECH_NOT U282 ( .A(n271), .Z(n267) );
  GTECH_OAI21 U283 ( .A(n310), .B(n311), .C(n312), .Z(n271) );
  GTECH_NOT U284 ( .A(n313), .Z(n272) );
  GTECH_NAND2 U285 ( .A(I_b[5]), .B(I_a[2]), .Z(n313) );
  GTECH_NOT U286 ( .A(n268), .Z(n270) );
  GTECH_NAND2 U287 ( .A(I_b[4]), .B(I_a[3]), .Z(n268) );
  GTECH_NOT U288 ( .A(n314), .Z(n276) );
  GTECH_NAND3 U289 ( .A(I_a[0]), .B(n315), .C(I_b[6]), .Z(n314) );
  GTECH_NOT U290 ( .A(n316), .Z(n315) );
  GTECH_NOT U291 ( .A(n260), .Z(n285) );
  GTECH_XNOR3 U292 ( .A(n280), .B(n282), .C(n277), .Z(n260) );
  GTECH_NOT U293 ( .A(n281), .Z(n277) );
  GTECH_OAI21 U294 ( .A(n317), .B(n318), .C(n319), .Z(n281) );
  GTECH_OAI21 U295 ( .A(n320), .B(n321), .C(n322), .Z(n319) );
  GTECH_NOT U296 ( .A(n323), .Z(n282) );
  GTECH_NAND2 U297 ( .A(I_b[3]), .B(I_a[4]), .Z(n323) );
  GTECH_NOT U298 ( .A(n278), .Z(n280) );
  GTECH_NAND2 U299 ( .A(I_a[5]), .B(I_b[2]), .Z(n278) );
  GTECH_NOT U300 ( .A(n324), .Z(n259) );
  GTECH_XNOR3 U301 ( .A(n286), .B(n287), .C(n290), .Z(n324) );
  GTECH_NOT U302 ( .A(n288), .Z(n290) );
  GTECH_OAI21 U303 ( .A(n325), .B(n326), .C(n327), .Z(n288) );
  GTECH_OAI21 U304 ( .A(n305), .B(n307), .C(n306), .Z(n327) );
  GTECH_NOT U305 ( .A(n328), .Z(n287) );
  GTECH_NAND2 U306 ( .A(I_a[6]), .B(I_b[1]), .Z(n328) );
  GTECH_NOT U307 ( .A(n291), .Z(n286) );
  GTECH_NAND2 U308 ( .A(I_a[7]), .B(I_b[0]), .Z(n291) );
  GTECH_XOR2 U309 ( .A(n329), .B(n330), .Z(N146) );
  GTECH_OA21 U310 ( .A(n300), .B(n301), .C(n302), .Z(n330) );
  GTECH_OAI21 U311 ( .A(n331), .B(n332), .C(n333), .Z(n302) );
  GTECH_XOR4 U312 ( .A(n298), .B(n297), .C(n299), .D(n296), .Z(n329) );
  GTECH_XOR2 U313 ( .A(n316), .B(n334), .Z(n296) );
  GTECH_AND2 U314 ( .A(I_b[6]), .B(I_a[0]), .Z(n334) );
  GTECH_XNOR3 U315 ( .A(n335), .B(n336), .C(n337), .Z(n316) );
  GTECH_NOT U316 ( .A(n312), .Z(n337) );
  GTECH_NAND3 U317 ( .A(I_b[4]), .B(I_a[1]), .C(n338), .Z(n312) );
  GTECH_NOT U318 ( .A(n311), .Z(n336) );
  GTECH_NAND2 U319 ( .A(I_b[5]), .B(I_a[1]), .Z(n311) );
  GTECH_NOT U320 ( .A(n310), .Z(n335) );
  GTECH_NAND2 U321 ( .A(I_b[4]), .B(I_a[2]), .Z(n310) );
  GTECH_XNOR3 U322 ( .A(n320), .B(n322), .C(n317), .Z(n299) );
  GTECH_NOT U323 ( .A(n321), .Z(n317) );
  GTECH_OAI21 U324 ( .A(n339), .B(n340), .C(n341), .Z(n321) );
  GTECH_OAI21 U325 ( .A(n342), .B(n343), .C(n344), .Z(n341) );
  GTECH_NOT U326 ( .A(n345), .Z(n322) );
  GTECH_NAND2 U327 ( .A(I_b[3]), .B(I_a[3]), .Z(n345) );
  GTECH_NOT U328 ( .A(n318), .Z(n320) );
  GTECH_NAND2 U329 ( .A(I_b[2]), .B(I_a[4]), .Z(n318) );
  GTECH_ADD_ABC U330 ( .A(n346), .B(n347), .C(n348), .COUT(n297) );
  GTECH_NOT U331 ( .A(n349), .Z(n348) );
  GTECH_XNOR3 U332 ( .A(n350), .B(n351), .C(n352), .Z(n347) );
  GTECH_NOT U333 ( .A(n353), .Z(n298) );
  GTECH_XNOR3 U334 ( .A(n305), .B(n306), .C(n325), .Z(n353) );
  GTECH_NOT U335 ( .A(n307), .Z(n325) );
  GTECH_OAI21 U336 ( .A(n354), .B(n355), .C(n356), .Z(n307) );
  GTECH_OAI21 U337 ( .A(n350), .B(n352), .C(n351), .Z(n356) );
  GTECH_NOT U338 ( .A(n357), .Z(n306) );
  GTECH_NAND2 U339 ( .A(I_a[5]), .B(I_b[1]), .Z(n357) );
  GTECH_NOT U340 ( .A(n326), .Z(n305) );
  GTECH_NAND2 U341 ( .A(I_a[6]), .B(I_b[0]), .Z(n326) );
  GTECH_XNOR3 U342 ( .A(n333), .B(n301), .C(n332), .Z(N145) );
  GTECH_NOT U343 ( .A(n300), .Z(n332) );
  GTECH_XOR2 U344 ( .A(n358), .B(n338), .Z(n300) );
  GTECH_NOT U345 ( .A(n359), .Z(n338) );
  GTECH_NAND2 U346 ( .A(I_b[5]), .B(I_a[0]), .Z(n359) );
  GTECH_NAND2 U347 ( .A(I_b[4]), .B(I_a[1]), .Z(n358) );
  GTECH_NOT U348 ( .A(n331), .Z(n301) );
  GTECH_XOR2 U349 ( .A(n360), .B(n346), .Z(n331) );
  GTECH_ADD_ABC U350 ( .A(n361), .B(n362), .C(n363), .COUT(n346) );
  GTECH_XNOR3 U351 ( .A(n364), .B(n365), .C(n366), .Z(n362) );
  GTECH_OA21 U352 ( .A(n367), .B(n368), .C(n369), .Z(n361) );
  GTECH_XOR4 U353 ( .A(n351), .B(n354), .C(n349), .D(n350), .Z(n360) );
  GTECH_NOT U354 ( .A(n355), .Z(n350) );
  GTECH_NAND2 U355 ( .A(I_a[5]), .B(I_b[0]), .Z(n355) );
  GTECH_XNOR3 U356 ( .A(n342), .B(n344), .C(n339), .Z(n349) );
  GTECH_NOT U357 ( .A(n343), .Z(n339) );
  GTECH_OAI21 U358 ( .A(n370), .B(n371), .C(n372), .Z(n343) );
  GTECH_NOT U359 ( .A(n373), .Z(n344) );
  GTECH_NAND2 U360 ( .A(I_b[3]), .B(I_a[2]), .Z(n373) );
  GTECH_NOT U361 ( .A(n340), .Z(n342) );
  GTECH_NAND2 U362 ( .A(I_b[2]), .B(I_a[3]), .Z(n340) );
  GTECH_NOT U363 ( .A(n352), .Z(n354) );
  GTECH_OAI21 U364 ( .A(n374), .B(n375), .C(n376), .Z(n352) );
  GTECH_OAI21 U365 ( .A(n364), .B(n366), .C(n365), .Z(n376) );
  GTECH_NOT U366 ( .A(n375), .Z(n364) );
  GTECH_NOT U367 ( .A(n377), .Z(n351) );
  GTECH_NAND2 U368 ( .A(I_a[4]), .B(I_b[1]), .Z(n377) );
  GTECH_NOT U369 ( .A(n378), .Z(n333) );
  GTECH_NAND3 U370 ( .A(I_a[0]), .B(n379), .C(I_b[4]), .Z(n378) );
  GTECH_XOR2 U371 ( .A(n380), .B(n379), .Z(N144) );
  GTECH_XOR2 U372 ( .A(n381), .B(n382), .Z(n379) );
  GTECH_OA21 U373 ( .A(n367), .B(n368), .C(n369), .Z(n382) );
  GTECH_OAI21 U374 ( .A(n383), .B(n384), .C(n385), .Z(n369) );
  GTECH_XOR4 U375 ( .A(n365), .B(n374), .C(n375), .D(n363), .Z(n381) );
  GTECH_XNOR3 U376 ( .A(n386), .B(n387), .C(n388), .Z(n363) );
  GTECH_NOT U377 ( .A(n372), .Z(n388) );
  GTECH_NAND3 U378 ( .A(I_b[2]), .B(I_a[1]), .C(n389), .Z(n372) );
  GTECH_NOT U379 ( .A(n371), .Z(n387) );
  GTECH_NAND2 U380 ( .A(I_b[3]), .B(I_a[1]), .Z(n371) );
  GTECH_NOT U381 ( .A(n370), .Z(n386) );
  GTECH_NAND2 U382 ( .A(I_b[2]), .B(I_a[2]), .Z(n370) );
  GTECH_NAND2 U383 ( .A(I_a[4]), .B(I_b[0]), .Z(n375) );
  GTECH_NOT U384 ( .A(n366), .Z(n374) );
  GTECH_OAI21 U385 ( .A(n390), .B(n391), .C(n392), .Z(n366) );
  GTECH_OAI21 U386 ( .A(n393), .B(n394), .C(n395), .Z(n392) );
  GTECH_NOT U387 ( .A(n396), .Z(n365) );
  GTECH_NAND2 U388 ( .A(I_a[3]), .B(I_b[1]), .Z(n396) );
  GTECH_AND2 U389 ( .A(I_b[4]), .B(I_a[0]), .Z(n380) );
  GTECH_XNOR3 U390 ( .A(n385), .B(n368), .C(n384), .Z(N143) );
  GTECH_NOT U391 ( .A(n367), .Z(n384) );
  GTECH_XOR2 U392 ( .A(n397), .B(n389), .Z(n367) );
  GTECH_NOT U393 ( .A(n398), .Z(n389) );
  GTECH_NAND2 U394 ( .A(I_b[3]), .B(I_a[0]), .Z(n398) );
  GTECH_NAND2 U395 ( .A(I_b[2]), .B(I_a[1]), .Z(n397) );
  GTECH_NOT U396 ( .A(n383), .Z(n368) );
  GTECH_XNOR3 U397 ( .A(n393), .B(n395), .C(n390), .Z(n383) );
  GTECH_NOT U398 ( .A(n394), .Z(n390) );
  GTECH_OAI21 U399 ( .A(n399), .B(n400), .C(n401), .Z(n394) );
  GTECH_NOT U400 ( .A(n402), .Z(n395) );
  GTECH_NAND2 U401 ( .A(I_b[1]), .B(I_a[2]), .Z(n402) );
  GTECH_NOT U402 ( .A(n391), .Z(n393) );
  GTECH_NAND2 U403 ( .A(I_b[0]), .B(I_a[3]), .Z(n391) );
  GTECH_NOT U404 ( .A(n403), .Z(n385) );
  GTECH_NAND3 U405 ( .A(I_a[0]), .B(n404), .C(I_b[2]), .Z(n403) );
  GTECH_XOR2 U406 ( .A(n405), .B(n404), .Z(N142) );
  GTECH_NOT U407 ( .A(n406), .Z(n404) );
  GTECH_XNOR3 U408 ( .A(n407), .B(n408), .C(n409), .Z(n406) );
  GTECH_NOT U409 ( .A(n401), .Z(n409) );
  GTECH_NAND3 U410 ( .A(n410), .B(I_b[0]), .C(I_a[1]), .Z(n401) );
  GTECH_NOT U411 ( .A(n399), .Z(n408) );
  GTECH_NAND2 U412 ( .A(I_a[1]), .B(I_b[1]), .Z(n399) );
  GTECH_NOT U413 ( .A(n400), .Z(n407) );
  GTECH_NAND2 U414 ( .A(I_b[0]), .B(I_a[2]), .Z(n400) );
  GTECH_AND2 U415 ( .A(I_b[2]), .B(I_a[0]), .Z(n405) );
  GTECH_XOR2 U416 ( .A(n410), .B(n411), .Z(N141) );
  GTECH_AND2 U417 ( .A(I_a[1]), .B(I_b[0]), .Z(n411) );
  GTECH_NOT U418 ( .A(n412), .Z(n410) );
  GTECH_NAND2 U419 ( .A(I_a[0]), .B(I_b[1]), .Z(n412) );
  GTECH_AND2 U420 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

