
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367;

  GTECH_MUX2 U131 ( .A(n270), .B(n271), .S(n272), .Z(sum[9]) );
  GTECH_XNOR2 U132 ( .A(n273), .B(n274), .Z(n271) );
  GTECH_XNOR2 U133 ( .A(n275), .B(n274), .Z(n270) );
  GTECH_OR_NOT U134 ( .A(n276), .B(n277), .Z(n274) );
  GTECH_NAND2 U135 ( .A(n278), .B(n279), .Z(sum[8]) );
  GTECH_AO21 U136 ( .A(n280), .B(n275), .C(n272), .Z(n279) );
  GTECH_MUX2 U137 ( .A(n281), .B(n282), .S(n283), .Z(sum[7]) );
  GTECH_XNOR2 U138 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_XOR2 U139 ( .A(n284), .B(n286), .Z(n281) );
  GTECH_OA21 U140 ( .A(n287), .B(n288), .C(n289), .Z(n286) );
  GTECH_XNOR2 U141 ( .A(a[7]), .B(b[7]), .Z(n284) );
  GTECH_MUX2 U142 ( .A(n290), .B(n291), .S(n283), .Z(sum[6]) );
  GTECH_XOR2 U143 ( .A(n292), .B(n293), .Z(n291) );
  GTECH_XOR2 U144 ( .A(n288), .B(n293), .Z(n290) );
  GTECH_NAND2 U145 ( .A(n294), .B(n289), .Z(n293) );
  GTECH_AOI21 U146 ( .A(n295), .B(n296), .C(n297), .Z(n288) );
  GTECH_MUX2 U147 ( .A(n298), .B(n299), .S(n300), .Z(sum[5]) );
  GTECH_OR_NOT U148 ( .A(n297), .B(n295), .Z(n300) );
  GTECH_AO21 U149 ( .A(n301), .B(n283), .C(n296), .Z(n299) );
  GTECH_OAI21 U150 ( .A(a[4]), .B(n283), .C(n302), .Z(n298) );
  GTECH_AO21 U151 ( .A(n283), .B(a[4]), .C(b[4]), .Z(n302) );
  GTECH_XNOR2 U152 ( .A(n283), .B(n303), .Z(sum[4]) );
  GTECH_MUX2 U153 ( .A(n304), .B(n305), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U154 ( .A(n306), .B(n307), .Z(n305) );
  GTECH_XOR2 U155 ( .A(n306), .B(n308), .Z(n304) );
  GTECH_OA21 U156 ( .A(n309), .B(n310), .C(n311), .Z(n308) );
  GTECH_XNOR2 U157 ( .A(a[3]), .B(b[3]), .Z(n306) );
  GTECH_MUX2 U158 ( .A(n312), .B(n313), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U159 ( .A(n314), .B(n315), .Z(n313) );
  GTECH_XNOR2 U160 ( .A(n310), .B(n314), .Z(n312) );
  GTECH_AND2 U161 ( .A(n316), .B(n311), .Z(n314) );
  GTECH_AOI21 U162 ( .A(n317), .B(n318), .C(n319), .Z(n310) );
  GTECH_MUX2 U163 ( .A(n320), .B(n321), .S(n322), .Z(sum[1]) );
  GTECH_OR_NOT U164 ( .A(n319), .B(n317), .Z(n322) );
  GTECH_AO21 U165 ( .A(n323), .B(cin), .C(n318), .Z(n321) );
  GTECH_OAI21 U166 ( .A(cin), .B(n318), .C(n323), .Z(n320) );
  GTECH_AND2 U167 ( .A(a[0]), .B(b[0]), .Z(n318) );
  GTECH_MUX2 U168 ( .A(n324), .B(n325), .S(n326), .Z(sum[15]) );
  GTECH_XOR2 U169 ( .A(n327), .B(n328), .Z(n325) );
  GTECH_AOI21 U170 ( .A(n329), .B(n330), .C(n331), .Z(n328) );
  GTECH_XNOR2 U171 ( .A(n327), .B(n332), .Z(n324) );
  GTECH_XNOR2 U172 ( .A(a[15]), .B(b[15]), .Z(n327) );
  GTECH_MUX2 U173 ( .A(n333), .B(n334), .S(n326), .Z(sum[14]) );
  GTECH_XNOR2 U174 ( .A(n330), .B(n335), .Z(n334) );
  GTECH_AO21 U175 ( .A(n336), .B(n337), .C(n338), .Z(n330) );
  GTECH_XNOR2 U176 ( .A(n335), .B(n339), .Z(n333) );
  GTECH_OR_NOT U177 ( .A(n331), .B(n329), .Z(n335) );
  GTECH_MUX2 U178 ( .A(n340), .B(n341), .S(n326), .Z(sum[13]) );
  GTECH_XOR2 U179 ( .A(n342), .B(n343), .Z(n341) );
  GTECH_XNOR2 U180 ( .A(n343), .B(n344), .Z(n340) );
  GTECH_OR_NOT U181 ( .A(n338), .B(n336), .Z(n343) );
  GTECH_NAND2 U182 ( .A(n345), .B(n346), .Z(sum[12]) );
  GTECH_AO21 U183 ( .A(n342), .B(n344), .C(n326), .Z(n346) );
  GTECH_MUX2 U184 ( .A(n347), .B(n348), .S(n272), .Z(sum[11]) );
  GTECH_XOR2 U185 ( .A(n349), .B(n350), .Z(n348) );
  GTECH_AOI21 U186 ( .A(n351), .B(n352), .C(n353), .Z(n350) );
  GTECH_XNOR2 U187 ( .A(n349), .B(n354), .Z(n347) );
  GTECH_XNOR2 U188 ( .A(a[11]), .B(b[11]), .Z(n349) );
  GTECH_MUX2 U189 ( .A(n355), .B(n356), .S(n272), .Z(sum[10]) );
  GTECH_XNOR2 U190 ( .A(n352), .B(n357), .Z(n356) );
  GTECH_AO21 U191 ( .A(n277), .B(n273), .C(n276), .Z(n352) );
  GTECH_NOT U192 ( .A(n280), .Z(n273) );
  GTECH_XNOR2 U193 ( .A(n358), .B(n357), .Z(n355) );
  GTECH_OR_NOT U194 ( .A(n353), .B(n351), .Z(n357) );
  GTECH_XOR2 U195 ( .A(cin), .B(n359), .Z(sum[0]) );
  GTECH_OAI21 U196 ( .A(n326), .B(n360), .C(n345), .Z(cout) );
  GTECH_NAND3 U197 ( .A(n342), .B(n344), .C(n326), .Z(n345) );
  GTECH_NOT U198 ( .A(n337), .Z(n342) );
  GTECH_AND2 U199 ( .A(b[12]), .B(a[12]), .Z(n337) );
  GTECH_AOI21 U200 ( .A(n332), .B(a[15]), .C(n361), .Z(n360) );
  GTECH_OA21 U201 ( .A(a[15]), .B(n332), .C(b[15]), .Z(n361) );
  GTECH_AO21 U202 ( .A(n339), .B(n329), .C(n331), .Z(n332) );
  GTECH_AND2 U203 ( .A(b[14]), .B(a[14]), .Z(n331) );
  GTECH_OR2 U204 ( .A(b[14]), .B(a[14]), .Z(n329) );
  GTECH_AO21 U205 ( .A(n336), .B(n344), .C(n338), .Z(n339) );
  GTECH_AND2 U206 ( .A(b[13]), .B(a[13]), .Z(n338) );
  GTECH_OR2 U207 ( .A(b[12]), .B(a[12]), .Z(n344) );
  GTECH_OR2 U208 ( .A(a[13]), .B(b[13]), .Z(n336) );
  GTECH_OA21 U209 ( .A(n362), .B(n272), .C(n278), .Z(n326) );
  GTECH_NAND3 U210 ( .A(n275), .B(n280), .C(n272), .Z(n278) );
  GTECH_NAND2 U211 ( .A(b[8]), .B(a[8]), .Z(n280) );
  GTECH_MUX2 U212 ( .A(n303), .B(n363), .S(n283), .Z(n272) );
  GTECH_MUX2 U213 ( .A(n359), .B(n364), .S(cin), .Z(n283) );
  GTECH_OA21 U214 ( .A(a[3]), .B(n307), .C(n365), .Z(n364) );
  GTECH_AO21 U215 ( .A(n307), .B(a[3]), .C(b[3]), .Z(n365) );
  GTECH_OAI21 U216 ( .A(n315), .B(n309), .C(n311), .Z(n307) );
  GTECH_NAND2 U217 ( .A(b[2]), .B(a[2]), .Z(n311) );
  GTECH_NOT U218 ( .A(n316), .Z(n309) );
  GTECH_OR2 U219 ( .A(b[2]), .B(a[2]), .Z(n316) );
  GTECH_AOI21 U220 ( .A(n323), .B(n317), .C(n319), .Z(n315) );
  GTECH_AND2 U221 ( .A(a[1]), .B(b[1]), .Z(n319) );
  GTECH_OR2 U222 ( .A(a[1]), .B(b[1]), .Z(n317) );
  GTECH_OR2 U223 ( .A(a[0]), .B(b[0]), .Z(n323) );
  GTECH_XOR2 U224 ( .A(a[0]), .B(b[0]), .Z(n359) );
  GTECH_OAI21 U225 ( .A(a[7]), .B(n285), .C(n366), .Z(n363) );
  GTECH_AO21 U226 ( .A(n285), .B(a[7]), .C(b[7]), .Z(n366) );
  GTECH_OAI21 U227 ( .A(n292), .B(n287), .C(n289), .Z(n285) );
  GTECH_NAND2 U228 ( .A(b[6]), .B(a[6]), .Z(n289) );
  GTECH_NOT U229 ( .A(n294), .Z(n287) );
  GTECH_OR2 U230 ( .A(b[6]), .B(a[6]), .Z(n294) );
  GTECH_AOI21 U231 ( .A(n301), .B(n295), .C(n297), .Z(n292) );
  GTECH_AND2 U232 ( .A(b[5]), .B(a[5]), .Z(n297) );
  GTECH_OR2 U233 ( .A(b[5]), .B(a[5]), .Z(n295) );
  GTECH_OR_NOT U234 ( .A(n296), .B(n301), .Z(n303) );
  GTECH_OR2 U235 ( .A(b[4]), .B(a[4]), .Z(n301) );
  GTECH_AND2 U236 ( .A(b[4]), .B(a[4]), .Z(n296) );
  GTECH_AOI21 U237 ( .A(n354), .B(a[11]), .C(n367), .Z(n362) );
  GTECH_OA21 U238 ( .A(a[11]), .B(n354), .C(b[11]), .Z(n367) );
  GTECH_AO21 U239 ( .A(n358), .B(n351), .C(n353), .Z(n354) );
  GTECH_AND2 U240 ( .A(b[10]), .B(a[10]), .Z(n353) );
  GTECH_OR2 U241 ( .A(b[10]), .B(a[10]), .Z(n351) );
  GTECH_AO21 U242 ( .A(n277), .B(n275), .C(n276), .Z(n358) );
  GTECH_AND2 U243 ( .A(b[9]), .B(a[9]), .Z(n276) );
  GTECH_OR2 U244 ( .A(b[8]), .B(a[8]), .Z(n275) );
  GTECH_OR2 U245 ( .A(b[9]), .B(a[9]), .Z(n277) );
endmodule

