
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n3, n4, n7, n8, n11, n12, n15, n16, n19, n20, n23, n24, n27, n28, n31,
         n32, n35, n36, n39, n40, n43, n44, n47, n48, n51, n52, n55, n56, n59,
         n60, n63, n64, n67, n68, n71, n72, n75, n76, n79, n80, n83, n84, n87,
         n88, n91, n92, n95, n96, n99, n100, n103, n104, n107, n108, n111,
         n112, n115, n116, n119, n120, n123, n124, n127, n128, n134, n133,
         n132, n137, n136, n135, n140, n139, n138, n143, n142, n141, n146,
         n145, n144, n149, n148, n147, n152, n151, n150, n153, n154, n158,
         n159, n160, n161, n162, n166, n165, n164, n163, n167, n168, n169,
         n173, n174, n175, n176, n177, n181, n180, n179, n178, n182, n183,
         n184, n188, n189, n190, n191, n192, n196, n195, n194, n193, n197,
         n198, n199, n203, n204, n205, n206, n207, n211, n210, n209, n208,
         n212, n215, n214, n213;
  wire   [131:129] n;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  GTECH_NOT first_I_0 ( .A(cin), .Z(n212) );
  SELECT_OP first_C17 ( .DATA1(n207), .DATA2(n206), .CONTROL1(n198), 
        .CONTROL2(n199), .Z(n213) );
  GTECH_BUF first_B_1 ( .A(n212), .Z(n199) );
  GTECH_BUF first_B_0 ( .A(cin), .Z(n198) );
  SELECT_OP first_C16 ( .DATA1({n208, n209, n210, n211}), .DATA2({n203, n204, 
        n205, n206}), .CONTROL1(n198), .CONTROL2(n199), .Z(sum[3:0]) );
  GTECH_NOT genblk1_1__my_adder_I_0 ( .A(n213), .Z(n197) );
  SELECT_OP genblk1_1__my_adder_C17 ( .DATA1(n192), .DATA2(n191), .CONTROL1(
        n183), .CONTROL2(n184), .Z(n214) );
  GTECH_BUF genblk1_1__my_adder_B_1 ( .A(n197), .Z(n184) );
  GTECH_BUF genblk1_1__my_adder_B_0 ( .A(n213), .Z(n183) );
  SELECT_OP genblk1_1__my_adder_C16 ( .DATA1({n193, n194, n195, n196}), 
        .DATA2({n188, n189, n190, n191}), .CONTROL1(n183), .CONTROL2(n184), 
        .Z(sum[7:4]) );
  GTECH_NOT genblk1_2__my_adder_I_0 ( .A(n214), .Z(n182) );
  SELECT_OP genblk1_2__my_adder_C17 ( .DATA1(n177), .DATA2(n176), .CONTROL1(
        n168), .CONTROL2(n169), .Z(n215) );
  GTECH_BUF genblk1_2__my_adder_B_1 ( .A(n182), .Z(n169) );
  GTECH_BUF genblk1_2__my_adder_B_0 ( .A(n214), .Z(n168) );
  SELECT_OP genblk1_2__my_adder_C16 ( .DATA1({n178, n179, n180, n181}), 
        .DATA2({n173, n174, n175, n176}), .CONTROL1(n168), .CONTROL2(n169), 
        .Z(sum[11:8]) );
  GTECH_NOT genblk1_3__my_adder_I_0 ( .A(n215), .Z(n167) );
  SELECT_OP genblk1_3__my_adder_C17 ( .DATA1(n162), .DATA2(n161), .CONTROL1(
        n153), .CONTROL2(n154), .Z(cout) );
  GTECH_BUF genblk1_3__my_adder_B_1 ( .A(n167), .Z(n154) );
  GTECH_BUF genblk1_3__my_adder_B_0 ( .A(n215), .Z(n153) );
  SELECT_OP genblk1_3__my_adder_C16 ( .DATA1({n163, n164, n165, n166}), 
        .DATA2({n158, n159, n160, n161}), .CONTROL1(n153), .CONTROL2(n154), 
        .Z(sum[15:12]) );
  GTECH_XOR2 first_adder0_first_C8 ( .A(a[0]), .B(b[0]) );
  GTECH_AND2 first_adder0_first_C7 ( .A(a[0]), .B(b[0]) );
  ADD_UNS_OP first_adder0_first_add_11_2 ( .A({n128, n127}), .B(1'b0), .Z({
        n152, n206}) );
  ADD_UNS_OP first_adder0_first_add_11 ( .A(a[0]), .B(b[0]), .Z({n128, n127})
         );
  GTECH_XOR2 first_adder0_genblk1_1__my_adder_C8 ( .A(a[1]), .B(b[1]) );
  GTECH_AND2 first_adder0_genblk1_1__my_adder_C7 ( .A(a[1]), .B(b[1]) );
  ADD_UNS_OP first_adder0_genblk1_1__my_adder_add_11_2 ( .A({n124, n123}), .B(
        n152), .Z({n151, n205}) );
  ADD_UNS_OP first_adder0_genblk1_1__my_adder_add_11 ( .A(a[1]), .B(b[1]), .Z(
        {n124, n123}) );
  GTECH_XOR2 first_adder0_genblk1_2__my_adder_C8 ( .A(a[2]), .B(b[2]) );
  GTECH_AND2 first_adder0_genblk1_2__my_adder_C7 ( .A(a[2]), .B(b[2]) );
  ADD_UNS_OP first_adder0_genblk1_2__my_adder_add_11_2 ( .A({n120, n119}), .B(
        n151), .Z({n150, n204}) );
  ADD_UNS_OP first_adder0_genblk1_2__my_adder_add_11 ( .A(a[2]), .B(b[2]), .Z(
        {n120, n119}) );
  GTECH_XOR2 first_adder0_genblk1_3__my_adder_C8 ( .A(a[3]), .B(b[3]) );
  GTECH_AND2 first_adder0_genblk1_3__my_adder_C7 ( .A(a[3]), .B(b[3]) );
  ADD_UNS_OP first_adder0_genblk1_3__my_adder_add_11_2 ( .A({n116, n115}), .B(
        n150), .Z({SYNOPSYS_UNCONNECTED__0, n203}) );
  ADD_UNS_OP first_adder0_genblk1_3__my_adder_add_11 ( .A(a[3]), .B(b[3]), .Z(
        {n116, n115}) );
  GTECH_XOR2 first_adder1_first_C8 ( .A(a[0]), .B(b[0]) );
  GTECH_AND2 first_adder1_first_C7 ( .A(a[0]), .B(b[0]) );
  ADD_UNS_OP first_adder1_first_add_11_2 ( .A({n112, n111}), .B(1'b1), .Z({
        n149, n211}) );
  ADD_UNS_OP first_adder1_first_add_11 ( .A(a[0]), .B(b[0]), .Z({n112, n111})
         );
  GTECH_XOR2 first_adder1_genblk1_1__my_adder_C8 ( .A(a[1]), .B(b[1]) );
  GTECH_AND2 first_adder1_genblk1_1__my_adder_C7 ( .A(a[1]), .B(b[1]) );
  ADD_UNS_OP first_adder1_genblk1_1__my_adder_add_11_2 ( .A({n108, n107}), .B(
        n149), .Z({n148, n210}) );
  ADD_UNS_OP first_adder1_genblk1_1__my_adder_add_11 ( .A(a[1]), .B(b[1]), .Z(
        {n108, n107}) );
  GTECH_XOR2 first_adder1_genblk1_2__my_adder_C8 ( .A(a[2]), .B(b[2]) );
  GTECH_AND2 first_adder1_genblk1_2__my_adder_C7 ( .A(a[2]), .B(b[2]) );
  ADD_UNS_OP first_adder1_genblk1_2__my_adder_add_11_2 ( .A({n104, n103}), .B(
        n148), .Z({n147, n209}) );
  ADD_UNS_OP first_adder1_genblk1_2__my_adder_add_11 ( .A(a[2]), .B(b[2]), .Z(
        {n104, n103}) );
  GTECH_XOR2 first_adder1_genblk1_3__my_adder_C8 ( .A(a[3]), .B(b[3]) );
  GTECH_AND2 first_adder1_genblk1_3__my_adder_C7 ( .A(a[3]), .B(b[3]) );
  ADD_UNS_OP first_adder1_genblk1_3__my_adder_add_11_2 ( .A({n100, n99}), .B(
        n147), .Z({n207, n208}) );
  ADD_UNS_OP first_adder1_genblk1_3__my_adder_add_11 ( .A(a[3]), .B(b[3]), .Z(
        {n100, n99}) );
  GTECH_XOR2 genblk1_1__my_adder_adder0_first_C8 ( .A(a[4]), .B(b[4]) );
  GTECH_AND2 genblk1_1__my_adder_adder0_first_C7 ( .A(a[4]), .B(b[4]) );
  ADD_UNS_OP genblk1_1__my_adder_adder0_first_add_11_2 ( .A({n96, n95}), .B(
        1'b0), .Z({n146, n191}) );
  ADD_UNS_OP genblk1_1__my_adder_adder0_first_add_11 ( .A(a[4]), .B(b[4]), .Z(
        {n96, n95}) );
  GTECH_XOR2 genblk1_1__my_adder_adder0_genblk1_1__my_adder_C8 ( .A(a[5]), .B(
        b[5]) );
  GTECH_AND2 genblk1_1__my_adder_adder0_genblk1_1__my_adder_C7 ( .A(a[5]), .B(
        b[5]) );
  ADD_UNS_OP genblk1_1__my_adder_adder0_genblk1_1__my_adder_add_11_2 ( .A({n92, 
        n91}), .B(n146), .Z({n145, n190}) );
  ADD_UNS_OP genblk1_1__my_adder_adder0_genblk1_1__my_adder_add_11 ( .A(a[5]), 
        .B(b[5]), .Z({n92, n91}) );
  GTECH_XOR2 genblk1_1__my_adder_adder0_genblk1_2__my_adder_C8 ( .A(a[6]), .B(
        b[6]) );
  GTECH_AND2 genblk1_1__my_adder_adder0_genblk1_2__my_adder_C7 ( .A(a[6]), .B(
        b[6]) );
  ADD_UNS_OP genblk1_1__my_adder_adder0_genblk1_2__my_adder_add_11_2 ( .A({n88, 
        n87}), .B(n145), .Z({n144, n189}) );
  ADD_UNS_OP genblk1_1__my_adder_adder0_genblk1_2__my_adder_add_11 ( .A(a[6]), 
        .B(b[6]), .Z({n88, n87}) );
  GTECH_XOR2 genblk1_1__my_adder_adder0_genblk1_3__my_adder_C8 ( .A(a[7]), .B(
        b[7]) );
  GTECH_AND2 genblk1_1__my_adder_adder0_genblk1_3__my_adder_C7 ( .A(a[7]), .B(
        b[7]) );
  ADD_UNS_OP genblk1_1__my_adder_adder0_genblk1_3__my_adder_add_11_2 ( .A({n84, 
        n83}), .B(n144), .Z({SYNOPSYS_UNCONNECTED__1, n188}) );
  ADD_UNS_OP genblk1_1__my_adder_adder0_genblk1_3__my_adder_add_11 ( .A(a[7]), 
        .B(b[7]), .Z({n84, n83}) );
  GTECH_XOR2 genblk1_1__my_adder_adder1_first_C8 ( .A(a[4]), .B(b[4]) );
  GTECH_AND2 genblk1_1__my_adder_adder1_first_C7 ( .A(a[4]), .B(b[4]) );
  ADD_UNS_OP genblk1_1__my_adder_adder1_first_add_11_2 ( .A({n80, n79}), .B(
        1'b1), .Z({n143, n196}) );
  ADD_UNS_OP genblk1_1__my_adder_adder1_first_add_11 ( .A(a[4]), .B(b[4]), .Z(
        {n80, n79}) );
  GTECH_XOR2 genblk1_1__my_adder_adder1_genblk1_1__my_adder_C8 ( .A(a[5]), .B(
        b[5]) );
  GTECH_AND2 genblk1_1__my_adder_adder1_genblk1_1__my_adder_C7 ( .A(a[5]), .B(
        b[5]) );
  ADD_UNS_OP genblk1_1__my_adder_adder1_genblk1_1__my_adder_add_11_2 ( .A({n76, 
        n75}), .B(n143), .Z({n142, n195}) );
  ADD_UNS_OP genblk1_1__my_adder_adder1_genblk1_1__my_adder_add_11 ( .A(a[5]), 
        .B(b[5]), .Z({n76, n75}) );
  GTECH_XOR2 genblk1_1__my_adder_adder1_genblk1_2__my_adder_C8 ( .A(a[6]), .B(
        b[6]) );
  GTECH_AND2 genblk1_1__my_adder_adder1_genblk1_2__my_adder_C7 ( .A(a[6]), .B(
        b[6]) );
  ADD_UNS_OP genblk1_1__my_adder_adder1_genblk1_2__my_adder_add_11_2 ( .A({n72, 
        n71}), .B(n142), .Z({n141, n194}) );
  ADD_UNS_OP genblk1_1__my_adder_adder1_genblk1_2__my_adder_add_11 ( .A(a[6]), 
        .B(b[6]), .Z({n72, n71}) );
  GTECH_XOR2 genblk1_1__my_adder_adder1_genblk1_3__my_adder_C8 ( .A(a[7]), .B(
        b[7]) );
  GTECH_AND2 genblk1_1__my_adder_adder1_genblk1_3__my_adder_C7 ( .A(a[7]), .B(
        b[7]) );
  ADD_UNS_OP genblk1_1__my_adder_adder1_genblk1_3__my_adder_add_11_2 ( .A({n68, 
        n67}), .B(n141), .Z({n192, n193}) );
  ADD_UNS_OP genblk1_1__my_adder_adder1_genblk1_3__my_adder_add_11 ( .A(a[7]), 
        .B(b[7]), .Z({n68, n67}) );
  GTECH_XOR2 genblk1_2__my_adder_adder0_first_C8 ( .A(a[8]), .B(b[8]) );
  GTECH_AND2 genblk1_2__my_adder_adder0_first_C7 ( .A(a[8]), .B(b[8]) );
  ADD_UNS_OP genblk1_2__my_adder_adder0_first_add_11_2 ( .A({n64, n63}), .B(
        1'b0), .Z({n140, n176}) );
  ADD_UNS_OP genblk1_2__my_adder_adder0_first_add_11 ( .A(a[8]), .B(b[8]), .Z(
        {n64, n63}) );
  GTECH_XOR2 genblk1_2__my_adder_adder0_genblk1_1__my_adder_C8 ( .A(a[9]), .B(
        b[9]) );
  GTECH_AND2 genblk1_2__my_adder_adder0_genblk1_1__my_adder_C7 ( .A(a[9]), .B(
        b[9]) );
  ADD_UNS_OP genblk1_2__my_adder_adder0_genblk1_1__my_adder_add_11_2 ( .A({n60, 
        n59}), .B(n140), .Z({n139, n175}) );
  ADD_UNS_OP genblk1_2__my_adder_adder0_genblk1_1__my_adder_add_11 ( .A(a[9]), 
        .B(b[9]), .Z({n60, n59}) );
  GTECH_XOR2 genblk1_2__my_adder_adder0_genblk1_2__my_adder_C8 ( .A(a[10]), 
        .B(b[10]) );
  GTECH_AND2 genblk1_2__my_adder_adder0_genblk1_2__my_adder_C7 ( .A(a[10]), 
        .B(b[10]) );
  ADD_UNS_OP genblk1_2__my_adder_adder0_genblk1_2__my_adder_add_11_2 ( .A({n56, 
        n55}), .B(n139), .Z({n138, n174}) );
  ADD_UNS_OP genblk1_2__my_adder_adder0_genblk1_2__my_adder_add_11 ( .A(a[10]), 
        .B(b[10]), .Z({n56, n55}) );
  GTECH_XOR2 genblk1_2__my_adder_adder0_genblk1_3__my_adder_C8 ( .A(a[11]), 
        .B(b[11]) );
  GTECH_AND2 genblk1_2__my_adder_adder0_genblk1_3__my_adder_C7 ( .A(a[11]), 
        .B(b[11]) );
  ADD_UNS_OP genblk1_2__my_adder_adder0_genblk1_3__my_adder_add_11_2 ( .A({n52, 
        n51}), .B(n138), .Z({SYNOPSYS_UNCONNECTED__2, n173}) );
  ADD_UNS_OP genblk1_2__my_adder_adder0_genblk1_3__my_adder_add_11 ( .A(a[11]), 
        .B(b[11]), .Z({n52, n51}) );
  GTECH_XOR2 genblk1_2__my_adder_adder1_first_C8 ( .A(a[8]), .B(b[8]) );
  GTECH_AND2 genblk1_2__my_adder_adder1_first_C7 ( .A(a[8]), .B(b[8]) );
  ADD_UNS_OP genblk1_2__my_adder_adder1_first_add_11_2 ( .A({n48, n47}), .B(
        1'b1), .Z({n137, n181}) );
  ADD_UNS_OP genblk1_2__my_adder_adder1_first_add_11 ( .A(a[8]), .B(b[8]), .Z(
        {n48, n47}) );
  GTECH_XOR2 genblk1_2__my_adder_adder1_genblk1_1__my_adder_C8 ( .A(a[9]), .B(
        b[9]) );
  GTECH_AND2 genblk1_2__my_adder_adder1_genblk1_1__my_adder_C7 ( .A(a[9]), .B(
        b[9]) );
  ADD_UNS_OP genblk1_2__my_adder_adder1_genblk1_1__my_adder_add_11_2 ( .A({n44, 
        n43}), .B(n137), .Z({n136, n180}) );
  ADD_UNS_OP genblk1_2__my_adder_adder1_genblk1_1__my_adder_add_11 ( .A(a[9]), 
        .B(b[9]), .Z({n44, n43}) );
  GTECH_XOR2 genblk1_2__my_adder_adder1_genblk1_2__my_adder_C8 ( .A(a[10]), 
        .B(b[10]) );
  GTECH_AND2 genblk1_2__my_adder_adder1_genblk1_2__my_adder_C7 ( .A(a[10]), 
        .B(b[10]) );
  ADD_UNS_OP genblk1_2__my_adder_adder1_genblk1_2__my_adder_add_11_2 ( .A({n40, 
        n39}), .B(n136), .Z({n135, n179}) );
  ADD_UNS_OP genblk1_2__my_adder_adder1_genblk1_2__my_adder_add_11 ( .A(a[10]), 
        .B(b[10]), .Z({n40, n39}) );
  GTECH_XOR2 genblk1_2__my_adder_adder1_genblk1_3__my_adder_C8 ( .A(a[11]), 
        .B(b[11]) );
  GTECH_AND2 genblk1_2__my_adder_adder1_genblk1_3__my_adder_C7 ( .A(a[11]), 
        .B(b[11]) );
  ADD_UNS_OP genblk1_2__my_adder_adder1_genblk1_3__my_adder_add_11_2 ( .A({n36, 
        n35}), .B(n135), .Z({n177, n178}) );
  ADD_UNS_OP genblk1_2__my_adder_adder1_genblk1_3__my_adder_add_11 ( .A(a[11]), 
        .B(b[11]), .Z({n36, n35}) );
  GTECH_XOR2 genblk1_3__my_adder_adder0_first_C8 ( .A(a[12]), .B(b[12]) );
  GTECH_AND2 genblk1_3__my_adder_adder0_first_C7 ( .A(a[12]), .B(b[12]) );
  ADD_UNS_OP genblk1_3__my_adder_adder0_first_add_11_2 ( .A({n32, n31}), .B(
        1'b0), .Z({n134, n161}) );
  ADD_UNS_OP genblk1_3__my_adder_adder0_first_add_11 ( .A(a[12]), .B(b[12]), 
        .Z({n32, n31}) );
  GTECH_XOR2 genblk1_3__my_adder_adder0_genblk1_1__my_adder_C8 ( .A(a[13]), 
        .B(b[13]) );
  GTECH_AND2 genblk1_3__my_adder_adder0_genblk1_1__my_adder_C7 ( .A(a[13]), 
        .B(b[13]) );
  ADD_UNS_OP genblk1_3__my_adder_adder0_genblk1_1__my_adder_add_11_2 ( .A({n28, 
        n27}), .B(n134), .Z({n133, n160}) );
  ADD_UNS_OP genblk1_3__my_adder_adder0_genblk1_1__my_adder_add_11 ( .A(a[13]), 
        .B(b[13]), .Z({n28, n27}) );
  GTECH_XOR2 genblk1_3__my_adder_adder0_genblk1_2__my_adder_C8 ( .A(a[14]), 
        .B(b[14]) );
  GTECH_AND2 genblk1_3__my_adder_adder0_genblk1_2__my_adder_C7 ( .A(a[14]), 
        .B(b[14]) );
  ADD_UNS_OP genblk1_3__my_adder_adder0_genblk1_2__my_adder_add_11_2 ( .A({n24, 
        n23}), .B(n133), .Z({n132, n159}) );
  ADD_UNS_OP genblk1_3__my_adder_adder0_genblk1_2__my_adder_add_11 ( .A(a[14]), 
        .B(b[14]), .Z({n24, n23}) );
  GTECH_XOR2 genblk1_3__my_adder_adder0_genblk1_3__my_adder_C8 ( .A(a[15]), 
        .B(b[15]) );
  GTECH_AND2 genblk1_3__my_adder_adder0_genblk1_3__my_adder_C7 ( .A(a[15]), 
        .B(b[15]) );
  ADD_UNS_OP genblk1_3__my_adder_adder0_genblk1_3__my_adder_add_11_2 ( .A({n20, 
        n19}), .B(n132), .Z({SYNOPSYS_UNCONNECTED__3, n158}) );
  ADD_UNS_OP genblk1_3__my_adder_adder0_genblk1_3__my_adder_add_11 ( .A(a[15]), 
        .B(b[15]), .Z({n20, n19}) );
  GTECH_XOR2 genblk1_3__my_adder_adder1_first_C8 ( .A(a[12]), .B(b[12]) );
  GTECH_AND2 genblk1_3__my_adder_adder1_first_C7 ( .A(a[12]), .B(b[12]) );
  ADD_UNS_OP genblk1_3__my_adder_adder1_first_add_11_2 ( .A({n16, n15}), .B(
        1'b1), .Z({n[131], n166}) );
  ADD_UNS_OP genblk1_3__my_adder_adder1_first_add_11 ( .A(a[12]), .B(b[12]), 
        .Z({n16, n15}) );
  GTECH_XOR2 genblk1_3__my_adder_adder1_genblk1_1__my_adder_C8 ( .A(a[13]), 
        .B(b[13]) );
  GTECH_AND2 genblk1_3__my_adder_adder1_genblk1_1__my_adder_C7 ( .A(a[13]), 
        .B(b[13]) );
  ADD_UNS_OP genblk1_3__my_adder_adder1_genblk1_1__my_adder_add_11_2 ( .A({n12, 
        n11}), .B(n[131]), .Z({n[130], n165}) );
  ADD_UNS_OP genblk1_3__my_adder_adder1_genblk1_1__my_adder_add_11 ( .A(a[13]), 
        .B(b[13]), .Z({n12, n11}) );
  GTECH_XOR2 genblk1_3__my_adder_adder1_genblk1_2__my_adder_C8 ( .A(a[14]), 
        .B(b[14]) );
  GTECH_AND2 genblk1_3__my_adder_adder1_genblk1_2__my_adder_C7 ( .A(a[14]), 
        .B(b[14]) );
  ADD_UNS_OP genblk1_3__my_adder_adder1_genblk1_2__my_adder_add_11_2 ( .A({n8, 
        n7}), .B(n[130]), .Z({n[129], n164}) );
  ADD_UNS_OP genblk1_3__my_adder_adder1_genblk1_2__my_adder_add_11 ( .A(a[14]), 
        .B(b[14]), .Z({n8, n7}) );
  GTECH_XOR2 genblk1_3__my_adder_adder1_genblk1_3__my_adder_C8 ( .A(a[15]), 
        .B(b[15]) );
  GTECH_AND2 genblk1_3__my_adder_adder1_genblk1_3__my_adder_C7 ( .A(a[15]), 
        .B(b[15]) );
  ADD_UNS_OP genblk1_3__my_adder_adder1_genblk1_3__my_adder_add_11_2 ( .A({n4, 
        n3}), .B(n[129]), .Z({n162, n163}) );
  ADD_UNS_OP genblk1_3__my_adder_adder1_genblk1_3__my_adder_add_11 ( .A(a[15]), 
        .B(b[15]), .Z({n4, n3}) );
endmodule

