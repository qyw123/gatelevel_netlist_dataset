
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131;

  GTECH_XOR2 U86 ( .A(n67), .B(n68), .Z(sum[9]) );
  GTECH_XOR2 U87 ( .A(n69), .B(n70), .Z(sum[8]) );
  GTECH_XNOR2 U88 ( .A(n71), .B(n72), .Z(sum[7]) );
  GTECH_AOI21 U89 ( .A(n73), .B(n74), .C(n75), .Z(n72) );
  GTECH_XOR2 U90 ( .A(n73), .B(n74), .Z(sum[6]) );
  GTECH_AO21 U91 ( .A(n76), .B(n77), .C(n78), .Z(n74) );
  GTECH_XOR2 U92 ( .A(n77), .B(n76), .Z(sum[5]) );
  GTECH_AO21 U93 ( .A(n79), .B(n80), .C(n81), .Z(n76) );
  GTECH_XOR2 U94 ( .A(n79), .B(n80), .Z(sum[4]) );
  GTECH_XNOR2 U95 ( .A(n82), .B(n83), .Z(sum[3]) );
  GTECH_AOI21 U96 ( .A(n84), .B(n85), .C(n86), .Z(n83) );
  GTECH_XOR2 U97 ( .A(n84), .B(n85), .Z(sum[2]) );
  GTECH_AO22 U98 ( .A(n87), .B(n88), .C(b[1]), .D(a[1]), .Z(n85) );
  GTECH_XOR2 U99 ( .A(n88), .B(n87), .Z(sum[1]) );
  GTECH_OR2 U100 ( .A(n89), .B(n90), .Z(n87) );
  GTECH_XNOR2 U101 ( .A(n91), .B(n92), .Z(sum[15]) );
  GTECH_AOI21 U102 ( .A(n93), .B(n94), .C(n95), .Z(n92) );
  GTECH_XOR2 U103 ( .A(n93), .B(n94), .Z(sum[14]) );
  GTECH_AO22 U104 ( .A(b[13]), .B(a[13]), .C(n96), .D(n97), .Z(n94) );
  GTECH_XOR2 U105 ( .A(n97), .B(n96), .Z(sum[13]) );
  GTECH_AO22 U106 ( .A(cout), .B(n98), .C(a[12]), .D(b[12]), .Z(n96) );
  GTECH_XOR2 U107 ( .A(n98), .B(cout), .Z(sum[12]) );
  GTECH_XNOR2 U108 ( .A(n99), .B(n100), .Z(sum[11]) );
  GTECH_AOI21 U109 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_XOR2 U110 ( .A(n101), .B(n102), .Z(sum[10]) );
  GTECH_OAI2N2 U111 ( .A(n68), .B(n67), .C(b[9]), .D(a[9]), .Z(n102) );
  GTECH_NOT U112 ( .A(n104), .Z(n67) );
  GTECH_AOI22 U113 ( .A(a[8]), .B(b[8]), .C(n70), .D(n69), .Z(n68) );
  GTECH_XNOR2 U114 ( .A(cin), .B(n105), .Z(sum[0]) );
  GTECH_AO21 U115 ( .A(n70), .B(n106), .C(n107), .Z(cout) );
  GTECH_AO21 U116 ( .A(n79), .B(n108), .C(n109), .Z(n70) );
  GTECH_AO21 U117 ( .A(n89), .B(n110), .C(n111), .Z(n79) );
  GTECH_AND2 U118 ( .A(cin), .B(n112), .Z(n89) );
  GTECH_AND4 U119 ( .A(n106), .B(n108), .C(n110), .D(n112), .Z(Pm) );
  GTECH_NOT U120 ( .A(n105), .Z(n112) );
  GTECH_OAI21 U121 ( .A(b[0]), .B(a[0]), .C(n113), .Z(n105) );
  GTECH_NOT U122 ( .A(n90), .Z(n113) );
  GTECH_AND4 U123 ( .A(n114), .B(n82), .C(n84), .D(n88), .Z(n110) );
  GTECH_AO21 U124 ( .A(n115), .B(n106), .C(n107), .Z(Gm) );
  GTECH_AO22 U125 ( .A(n116), .B(n91), .C(b[15]), .D(a[15]), .Z(n107) );
  GTECH_AO21 U126 ( .A(n93), .B(n117), .C(n95), .Z(n116) );
  GTECH_AND2 U127 ( .A(a[14]), .B(b[14]), .Z(n95) );
  GTECH_AO21 U128 ( .A(b[13]), .B(a[13]), .C(n118), .Z(n117) );
  GTECH_AND3 U129 ( .A(a[12]), .B(n97), .C(b[12]), .Z(n118) );
  GTECH_AND4 U130 ( .A(n98), .B(n91), .C(n93), .D(n97), .Z(n106) );
  GTECH_XOR2 U131 ( .A(a[13]), .B(b[13]), .Z(n97) );
  GTECH_XOR2 U132 ( .A(a[14]), .B(b[14]), .Z(n93) );
  GTECH_XOR2 U133 ( .A(a[15]), .B(b[15]), .Z(n91) );
  GTECH_XOR2 U134 ( .A(a[12]), .B(b[12]), .Z(n98) );
  GTECH_AO21 U135 ( .A(n108), .B(n111), .C(n109), .Z(n115) );
  GTECH_AO22 U136 ( .A(n119), .B(n99), .C(b[11]), .D(a[11]), .Z(n109) );
  GTECH_AO21 U137 ( .A(n101), .B(n120), .C(n103), .Z(n119) );
  GTECH_AND2 U138 ( .A(a[10]), .B(b[10]), .Z(n103) );
  GTECH_AO21 U139 ( .A(b[9]), .B(a[9]), .C(n121), .Z(n120) );
  GTECH_AND3 U140 ( .A(a[8]), .B(n104), .C(b[8]), .Z(n121) );
  GTECH_NOT U141 ( .A(n122), .Z(n111) );
  GTECH_AOI222 U142 ( .A(a[7]), .B(b[7]), .C(n114), .D(n123), .E(n71), .F(n124), .Z(n122) );
  GTECH_AO21 U143 ( .A(n125), .B(n73), .C(n75), .Z(n124) );
  GTECH_AO21 U144 ( .A(n81), .B(n77), .C(n78), .Z(n125) );
  GTECH_AND2 U145 ( .A(a[5]), .B(b[5]), .Z(n78) );
  GTECH_AO22 U146 ( .A(n126), .B(n82), .C(b[3]), .D(a[3]), .Z(n123) );
  GTECH_XOR2 U147 ( .A(a[3]), .B(b[3]), .Z(n82) );
  GTECH_AO21 U148 ( .A(n84), .B(n127), .C(n86), .Z(n126) );
  GTECH_AND2 U149 ( .A(a[2]), .B(b[2]), .Z(n86) );
  GTECH_AO22 U150 ( .A(b[1]), .B(a[1]), .C(n88), .D(n90), .Z(n127) );
  GTECH_AND2 U151 ( .A(b[0]), .B(a[0]), .Z(n90) );
  GTECH_XOR2 U152 ( .A(a[1]), .B(b[1]), .Z(n88) );
  GTECH_XOR2 U153 ( .A(a[2]), .B(b[2]), .Z(n84) );
  GTECH_AND4 U154 ( .A(n73), .B(n80), .C(n71), .D(n77), .Z(n114) );
  GTECH_XOR2 U155 ( .A(a[5]), .B(b[5]), .Z(n77) );
  GTECH_XOR2 U156 ( .A(a[7]), .B(b[7]), .Z(n71) );
  GTECH_AOI21 U157 ( .A(n128), .B(n129), .C(n81), .Z(n80) );
  GTECH_AND2 U158 ( .A(b[4]), .B(a[4]), .Z(n81) );
  GTECH_NOT U159 ( .A(a[4]), .Z(n129) );
  GTECH_NOT U160 ( .A(b[4]), .Z(n128) );
  GTECH_AOI21 U161 ( .A(n130), .B(n131), .C(n75), .Z(n73) );
  GTECH_AND2 U162 ( .A(b[6]), .B(a[6]), .Z(n75) );
  GTECH_NOT U163 ( .A(a[6]), .Z(n131) );
  GTECH_NOT U164 ( .A(b[6]), .Z(n130) );
  GTECH_AND4 U165 ( .A(n69), .B(n99), .C(n101), .D(n104), .Z(n108) );
  GTECH_XOR2 U166 ( .A(a[9]), .B(b[9]), .Z(n104) );
  GTECH_XOR2 U167 ( .A(a[10]), .B(b[10]), .Z(n101) );
  GTECH_XOR2 U168 ( .A(a[11]), .B(b[11]), .Z(n99) );
  GTECH_XOR2 U169 ( .A(a[8]), .B(b[8]), .Z(n69) );
endmodule

