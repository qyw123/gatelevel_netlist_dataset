
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142;

  GTECH_XOR2 U94 ( .A(n75), .B(n76), .Z(sum[9]) );
  GTECH_XOR2 U95 ( .A(n77), .B(n78), .Z(sum[8]) );
  GTECH_NOT U96 ( .A(n79), .Z(sum[7]) );
  GTECH_XOR2 U97 ( .A(n80), .B(n81), .Z(n79) );
  GTECH_AOI21 U98 ( .A(n82), .B(n83), .C(n84), .Z(n81) );
  GTECH_XOR2 U99 ( .A(n83), .B(n82), .Z(sum[6]) );
  GTECH_AO21 U100 ( .A(n85), .B(n86), .C(n87), .Z(n82) );
  GTECH_XOR2 U101 ( .A(n86), .B(n85), .Z(sum[5]) );
  GTECH_AO22 U102 ( .A(a[4]), .B(b[4]), .C(n88), .D(n89), .Z(n85) );
  GTECH_XOR2 U103 ( .A(n89), .B(n88), .Z(sum[4]) );
  GTECH_XOR2 U104 ( .A(n90), .B(n91), .Z(sum[3]) );
  GTECH_AOI21 U105 ( .A(n92), .B(n93), .C(n94), .Z(n91) );
  GTECH_XOR2 U106 ( .A(n93), .B(n92), .Z(sum[2]) );
  GTECH_AO21 U107 ( .A(n95), .B(n96), .C(n97), .Z(n92) );
  GTECH_XOR2 U108 ( .A(n96), .B(n95), .Z(sum[1]) );
  GTECH_OR_NOT U109 ( .A(n98), .B(n99), .Z(n95) );
  GTECH_XOR2 U110 ( .A(n100), .B(n101), .Z(sum[15]) );
  GTECH_AOI21 U111 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  GTECH_NOT U112 ( .A(n105), .Z(n100) );
  GTECH_XOR2 U113 ( .A(n103), .B(n102), .Z(sum[14]) );
  GTECH_AO21 U114 ( .A(n106), .B(n107), .C(n108), .Z(n102) );
  GTECH_XOR2 U115 ( .A(n107), .B(n106), .Z(sum[13]) );
  GTECH_AO22 U116 ( .A(a[12]), .B(b[12]), .C(cout), .D(n109), .Z(n106) );
  GTECH_XOR2 U117 ( .A(n109), .B(cout), .Z(sum[12]) );
  GTECH_XOR2 U118 ( .A(n110), .B(n111), .Z(sum[11]) );
  GTECH_AOI21 U119 ( .A(n112), .B(n113), .C(n114), .Z(n111) );
  GTECH_XOR2 U120 ( .A(n113), .B(n112), .Z(sum[10]) );
  GTECH_AO21 U121 ( .A(n76), .B(n75), .C(n115), .Z(n112) );
  GTECH_AO21 U122 ( .A(n78), .B(n77), .C(n116), .Z(n76) );
  GTECH_NOT U123 ( .A(n117), .Z(n78) );
  GTECH_XOR2 U124 ( .A(cin), .B(n118), .Z(sum[0]) );
  GTECH_OAI21 U125 ( .A(n117), .B(n119), .C(n120), .Z(cout) );
  GTECH_OA21 U126 ( .A(n121), .B(n122), .C(n123), .Z(n117) );
  GTECH_NOT U127 ( .A(n88), .Z(n121) );
  GTECH_OAI21 U128 ( .A(n99), .B(n124), .C(n125), .Z(n88) );
  GTECH_OR_NOT U129 ( .A(n126), .B(cin), .Z(n99) );
  GTECH_NOR4 U130 ( .A(n126), .B(n124), .C(n122), .D(n119), .Z(Pm) );
  GTECH_NAND4 U131 ( .A(n127), .B(n128), .C(n93), .D(n96), .Z(n124) );
  GTECH_NOT U132 ( .A(n118), .Z(n126) );
  GTECH_XOR2 U133 ( .A(a[0]), .B(b[0]), .Z(n118) );
  GTECH_OAI21 U134 ( .A(n129), .B(n119), .C(n120), .Z(Gm) );
  GTECH_AOI21 U135 ( .A(b[15]), .B(a[15]), .C(n130), .Z(n120) );
  GTECH_OA21 U136 ( .A(n104), .B(n131), .C(n105), .Z(n130) );
  GTECH_OA21 U137 ( .A(n108), .B(n132), .C(n103), .Z(n131) );
  GTECH_AND3 U138 ( .A(a[12]), .B(n107), .C(b[12]), .Z(n132) );
  GTECH_AND2 U139 ( .A(b[13]), .B(a[13]), .Z(n108) );
  GTECH_AND2 U140 ( .A(a[14]), .B(b[14]), .Z(n104) );
  GTECH_NAND4 U141 ( .A(n109), .B(n105), .C(n103), .D(n107), .Z(n119) );
  GTECH_XOR2 U142 ( .A(a[13]), .B(b[13]), .Z(n107) );
  GTECH_XOR2 U143 ( .A(a[14]), .B(b[14]), .Z(n103) );
  GTECH_XOR2 U144 ( .A(a[15]), .B(b[15]), .Z(n105) );
  GTECH_XOR2 U145 ( .A(a[12]), .B(b[12]), .Z(n109) );
  GTECH_OA21 U146 ( .A(n125), .B(n122), .C(n123), .Z(n129) );
  GTECH_AOI2N2 U147 ( .A(b[11]), .B(a[11]), .C(n133), .D(n110), .Z(n123) );
  GTECH_NOT U148 ( .A(n134), .Z(n110) );
  GTECH_AOI21 U149 ( .A(n135), .B(n113), .C(n114), .Z(n133) );
  GTECH_AND2 U150 ( .A(a[10]), .B(b[10]), .Z(n114) );
  GTECH_AO21 U151 ( .A(n75), .B(n116), .C(n115), .Z(n135) );
  GTECH_AND2 U152 ( .A(a[9]), .B(b[9]), .Z(n115) );
  GTECH_AND2 U153 ( .A(b[8]), .B(a[8]), .Z(n116) );
  GTECH_NAND4 U154 ( .A(n77), .B(n134), .C(n113), .D(n75), .Z(n122) );
  GTECH_XOR2 U155 ( .A(a[9]), .B(b[9]), .Z(n75) );
  GTECH_XOR2 U156 ( .A(a[10]), .B(b[10]), .Z(n113) );
  GTECH_XOR2 U157 ( .A(a[11]), .B(b[11]), .Z(n134) );
  GTECH_XOR2 U158 ( .A(a[8]), .B(b[8]), .Z(n77) );
  GTECH_AOI222 U159 ( .A(a[7]), .B(b[7]), .C(n80), .D(n136), .E(n127), .F(n137), .Z(n125) );
  GTECH_OAI2N2 U160 ( .A(n138), .B(n90), .C(b[3]), .D(a[3]), .Z(n137) );
  GTECH_NOT U161 ( .A(n128), .Z(n90) );
  GTECH_XOR2 U162 ( .A(a[3]), .B(b[3]), .Z(n128) );
  GTECH_AOI21 U163 ( .A(n139), .B(n93), .C(n94), .Z(n138) );
  GTECH_AND2 U164 ( .A(a[2]), .B(b[2]), .Z(n94) );
  GTECH_XOR2 U165 ( .A(a[2]), .B(b[2]), .Z(n93) );
  GTECH_AO21 U166 ( .A(n96), .B(n98), .C(n97), .Z(n139) );
  GTECH_AND2 U167 ( .A(a[1]), .B(b[1]), .Z(n97) );
  GTECH_AND2 U168 ( .A(b[0]), .B(a[0]), .Z(n98) );
  GTECH_XOR2 U169 ( .A(a[1]), .B(b[1]), .Z(n96) );
  GTECH_NOT U170 ( .A(n140), .Z(n127) );
  GTECH_NAND4 U171 ( .A(n89), .B(n80), .C(n83), .D(n86), .Z(n140) );
  GTECH_XOR2 U172 ( .A(a[4]), .B(b[4]), .Z(n89) );
  GTECH_OR_NOT U173 ( .A(n84), .B(n141), .Z(n136) );
  GTECH_OAI21 U174 ( .A(n142), .B(n87), .C(n83), .Z(n141) );
  GTECH_XOR2 U175 ( .A(a[6]), .B(b[6]), .Z(n83) );
  GTECH_AND2 U176 ( .A(a[5]), .B(b[5]), .Z(n87) );
  GTECH_AND3 U177 ( .A(a[4]), .B(n86), .C(b[4]), .Z(n142) );
  GTECH_XOR2 U178 ( .A(a[5]), .B(b[5]), .Z(n86) );
  GTECH_AND2 U179 ( .A(a[6]), .B(b[6]), .Z(n84) );
  GTECH_XOR2 U180 ( .A(a[7]), .B(b[7]), .Z(n80) );
endmodule

