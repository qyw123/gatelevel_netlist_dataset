
module clock_12h ( clk, reset, ena, pm, hh, mm, ss );
  output [7:0] hh;
  output [7:0] mm;
  output [7:0] ss;
  input clk, reset, ena;
  output pm;
  wire   N22, N23, N24, N25, N26, N39, N40, N41, N42, N43, N55, N56, N57, N58,
         N59, N71, N72, N73, N74, N75, N88, N89, N90, N91, N92, N110, N112,
         N114, N115, N116, N121, N122, n3, n4, n5, n6, n7, n8, n9, n78, n103,
         n104, n105, n106, n107, n108, n109, n110, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195;

  GTECH_FJK1S ss_ones_reg_0_ ( .J(n78), .K(n78), .TI(N22), .TE(N25), .CP(clk), 
        .Q(ss[0]) );
  GTECH_FJK1S ss_ones_reg_3_ ( .J(n78), .K(n78), .TI(N26), .TE(N25), .CP(clk), 
        .Q(ss[3]) );
  GTECH_FJK1S ss_ones_reg_1_ ( .J(n78), .K(n78), .TI(N23), .TE(N25), .CP(clk), 
        .Q(ss[1]) );
  GTECH_FJK1S ss_ones_reg_2_ ( .J(n78), .K(n78), .TI(N24), .TE(N25), .CP(clk), 
        .Q(ss[2]) );
  GTECH_FJK1S ss_tens_reg_0_ ( .J(n78), .K(n78), .TI(N39), .TE(N42), .CP(clk), 
        .Q(ss[4]) );
  GTECH_FJK1S ss_tens_reg_3_ ( .J(n78), .K(n78), .TI(N43), .TE(N42), .CP(clk), 
        .Q(ss[7]) );
  GTECH_FJK1S ss_tens_reg_1_ ( .J(n78), .K(n78), .TI(N40), .TE(N42), .CP(clk), 
        .Q(ss[5]) );
  GTECH_FJK1S ss_tens_reg_2_ ( .J(n78), .K(n78), .TI(N41), .TE(N42), .CP(clk), 
        .Q(ss[6]) );
  GTECH_FJK1S mm_ones_reg_0_ ( .J(n78), .K(n78), .TI(N55), .TE(N58), .CP(clk), 
        .Q(mm[0]), .QN(n3) );
  GTECH_FJK1S mm_ones_reg_3_ ( .J(n78), .K(n78), .TI(N59), .TE(N58), .CP(clk), 
        .Q(mm[3]), .QN(n108) );
  GTECH_FJK1S mm_ones_reg_1_ ( .J(n78), .K(n78), .TI(N56), .TE(N58), .CP(clk), 
        .Q(mm[1]), .QN(n110) );
  GTECH_FJK1S mm_ones_reg_2_ ( .J(n78), .K(n78), .TI(N57), .TE(N58), .CP(clk), 
        .Q(mm[2]), .QN(n109) );
  GTECH_FJK1S mm_tens_reg_0_ ( .J(n78), .K(n78), .TI(N71), .TE(N74), .CP(clk), 
        .Q(mm[4]), .QN(n4) );
  GTECH_FJK1S mm_tens_reg_3_ ( .J(n78), .K(n78), .TI(N75), .TE(N74), .CP(clk), 
        .Q(mm[7]), .QN(n105) );
  GTECH_FJK1S mm_tens_reg_1_ ( .J(n78), .K(n78), .TI(N72), .TE(N74), .CP(clk), 
        .Q(mm[5]), .QN(n107) );
  GTECH_FJK1S mm_tens_reg_2_ ( .J(n78), .K(n78), .TI(N73), .TE(N74), .CP(clk), 
        .Q(mm[6]), .QN(n106) );
  GTECH_FJK1S hh_tens_reg_0_ ( .J(n78), .K(n78), .TI(N110), .TE(N115), .CP(clk), .Q(hh[4]), .QN(n5) );
  GTECH_FJK1S hh_tens_reg_2_ ( .J(n78), .K(n78), .TI(N114), .TE(N115), .CP(clk), .Q(hh[6]), .QN(n6) );
  GTECH_FJK1S hh_tens_reg_3_ ( .J(n78), .K(n78), .TI(N116), .TE(N115), .CP(clk), .Q(hh[7]), .QN(n7) );
  GTECH_FJK1S hh_ones_reg_0_ ( .J(n78), .K(n78), .TI(N88), .TE(N91), .CP(clk), 
        .Q(hh[0]), .QN(n103) );
  GTECH_FJK1S hh_ones_reg_1_ ( .J(n78), .K(n78), .TI(N89), .TE(N91), .CP(clk), 
        .Q(hh[1]), .QN(n104) );
  GTECH_FJK1S hh_ones_reg_2_ ( .J(n78), .K(n78), .TI(N90), .TE(N91), .CP(clk), 
        .Q(hh[2]), .QN(n118) );
  GTECH_FJK1S hh_ones_reg_3_ ( .J(n78), .K(n78), .TI(N92), .TE(N91), .CP(clk), 
        .Q(hh[3]), .QN(n8) );
  GTECH_FJK1S hh_tens_reg_1_ ( .J(n78), .K(n78), .TI(N112), .TE(N115), .CP(clk), .Q(hh[5]), .QN(n9) );
  GTECH_FJK1S pm_temp_reg ( .J(n78), .K(n78), .TI(N122), .TE(N121), .CP(clk), 
        .Q(pm) );
  GTECH_ZERO U127 ( .Z(n78) );
  GTECH_AND_NOT U128 ( .A(n119), .B(n120), .Z(N92) );
  GTECH_XOR2 U129 ( .A(n121), .B(n8), .Z(n119) );
  GTECH_OR2 U130 ( .A(n118), .B(n122), .Z(n121) );
  GTECH_NAND2 U131 ( .A(n123), .B(n124), .Z(N91) );
  GTECH_AND_NOT U132 ( .A(n125), .B(n120), .Z(N90) );
  GTECH_XOR2 U133 ( .A(n122), .B(n118), .Z(n125) );
  GTECH_NAND2 U134 ( .A(n126), .B(n127), .Z(n122) );
  GTECH_OAI21 U135 ( .A(n128), .B(n120), .C(n123), .Z(N89) );
  GTECH_XOR2 U136 ( .A(n127), .B(n104), .Z(n128) );
  GTECH_OAI22 U137 ( .A(n124), .B(n129), .C(n127), .D(n120), .Z(N88) );
  GTECH_NAND3 U138 ( .A(n130), .B(n129), .C(n131), .Z(n120) );
  GTECH_AND_NOT U139 ( .A(n132), .B(n133), .Z(N75) );
  GTECH_MUX2 U140 ( .A(n134), .B(n135), .S(n105), .Z(n132) );
  GTECH_AND_NOT U141 ( .A(n136), .B(n4), .Z(n135) );
  GTECH_OR2 U142 ( .A(n106), .B(n137), .Z(n134) );
  GTECH_AND_NOT U143 ( .A(n138), .B(n133), .Z(N73) );
  GTECH_XOR2 U144 ( .A(n137), .B(n106), .Z(n138) );
  GTECH_AND_NOT U145 ( .A(n139), .B(n133), .Z(N72) );
  GTECH_OA21 U146 ( .A(n140), .B(n141), .C(n137), .Z(n139) );
  GTECH_NAND2 U147 ( .A(n140), .B(n141), .Z(n137) );
  GTECH_NOT U148 ( .A(n107), .Z(n140) );
  GTECH_AND_NOT U149 ( .A(n4), .B(n133), .Z(N71) );
  GTECH_NAND3 U150 ( .A(n142), .B(n123), .C(n143), .Z(n133) );
  GTECH_AND_NOT U151 ( .A(n144), .B(n145), .Z(N59) );
  GTECH_XOR2 U152 ( .A(n146), .B(n108), .Z(n144) );
  GTECH_OR2 U153 ( .A(n109), .B(n147), .Z(n146) );
  GTECH_AND_NOT U154 ( .A(n148), .B(n145), .Z(N57) );
  GTECH_XOR2 U155 ( .A(n147), .B(n109), .Z(n148) );
  GTECH_AND_NOT U156 ( .A(n149), .B(n145), .Z(N56) );
  GTECH_OA21 U157 ( .A(n150), .B(n151), .C(n147), .Z(n149) );
  GTECH_NAND2 U158 ( .A(n150), .B(n151), .Z(n147) );
  GTECH_NOT U159 ( .A(n110), .Z(n150) );
  GTECH_AND_NOT U160 ( .A(n3), .B(n145), .Z(N55) );
  GTECH_NAND2 U161 ( .A(n152), .B(n153), .Z(n145) );
  GTECH_NOT U162 ( .A(N74), .Z(n153) );
  GTECH_NAND2 U163 ( .A(n123), .B(n154), .Z(N74) );
  GTECH_NOR2 U164 ( .A(n155), .B(n156), .Z(N43) );
  GTECH_MUX2 U165 ( .A(n157), .B(n158), .S(ss[7]), .Z(n156) );
  GTECH_AND_NOT U166 ( .A(ss[6]), .B(n159), .Z(n158) );
  GTECH_NAND2 U167 ( .A(ss[6]), .B(ss[4]), .Z(n157) );
  GTECH_AND_NOT U168 ( .A(n160), .B(n161), .Z(N41) );
  GTECH_XOR2 U169 ( .A(n159), .B(ss[6]), .Z(n161) );
  GTECH_AND_NOT U170 ( .A(n162), .B(n155), .Z(N40) );
  GTECH_OA21 U171 ( .A(ss[4]), .B(ss[5]), .C(n159), .Z(n162) );
  GTECH_NAND2 U172 ( .A(ss[5]), .B(ss[4]), .Z(n159) );
  GTECH_AND_NOT U173 ( .A(n160), .B(ss[4]), .Z(N39) );
  GTECH_NOT U174 ( .A(n155), .Z(n160) );
  GTECH_NAND2 U175 ( .A(n163), .B(n164), .Z(n155) );
  GTECH_NOT U176 ( .A(N58), .Z(n164) );
  GTECH_NAND2 U177 ( .A(n123), .B(n165), .Z(N58) );
  GTECH_AND_NOT U178 ( .A(n166), .B(n167), .Z(N26) );
  GTECH_XNOR2 U179 ( .A(n168), .B(ss[3]), .Z(n167) );
  GTECH_AND_NOT U180 ( .A(ss[2]), .B(n169), .Z(n168) );
  GTECH_NAND2 U181 ( .A(n123), .B(n170), .Z(N25) );
  GTECH_NOT U182 ( .A(ena), .Z(n170) );
  GTECH_AND_NOT U183 ( .A(n166), .B(n171), .Z(N24) );
  GTECH_XOR2 U184 ( .A(n169), .B(ss[2]), .Z(n171) );
  GTECH_AND_NOT U185 ( .A(n172), .B(n173), .Z(N23) );
  GTECH_OA21 U186 ( .A(ss[0]), .B(ss[1]), .C(n169), .Z(n172) );
  GTECH_NAND2 U187 ( .A(ss[1]), .B(ss[0]), .Z(n169) );
  GTECH_AND_NOT U188 ( .A(n166), .B(ss[0]), .Z(N22) );
  GTECH_NOT U189 ( .A(n173), .Z(n166) );
  GTECH_NAND2 U190 ( .A(ena), .B(n174), .Z(n173) );
  GTECH_NOT U191 ( .A(N42), .Z(n174) );
  GTECH_NAND2 U192 ( .A(n123), .B(n175), .Z(N42) );
  GTECH_AND_NOT U193 ( .A(n176), .B(pm), .Z(N122) );
  GTECH_NOT U194 ( .A(n177), .Z(n176) );
  GTECH_NAND2 U195 ( .A(n123), .B(n177), .Z(N121) );
  GTECH_NAND4 U196 ( .A(n131), .B(n104), .C(n178), .D(n127), .Z(n177) );
  GTECH_AND_NOT U197 ( .A(n179), .B(n180), .Z(N116) );
  GTECH_XOR2 U198 ( .A(n181), .B(n7), .Z(n179) );
  GTECH_OR2 U199 ( .A(n6), .B(n182), .Z(n181) );
  GTECH_NAND3 U200 ( .A(n129), .B(n123), .C(n130), .Z(N115) );
  GTECH_NAND4 U201 ( .A(n103), .B(n178), .C(n183), .D(n126), .Z(n129) );
  GTECH_NOT U202 ( .A(n104), .Z(n126) );
  GTECH_AND3 U203 ( .A(n8), .B(n7), .C(n184), .Z(n178) );
  GTECH_AND4 U204 ( .A(n185), .B(n6), .C(n118), .D(n9), .Z(n184) );
  GTECH_AND_NOT U205 ( .A(n186), .B(n180), .Z(N114) );
  GTECH_XOR2 U206 ( .A(n182), .B(n6), .Z(n186) );
  GTECH_AND_NOT U207 ( .A(n187), .B(n180), .Z(N112) );
  GTECH_OA21 U208 ( .A(n188), .B(n185), .C(n182), .Z(n187) );
  GTECH_NAND2 U209 ( .A(n185), .B(n188), .Z(n182) );
  GTECH_NOT U210 ( .A(n9), .Z(n188) );
  GTECH_OAI21 U211 ( .A(n180), .B(n185), .C(n123), .Z(N110) );
  GTECH_NOT U212 ( .A(n5), .Z(n185) );
  GTECH_NAND2 U213 ( .A(n189), .B(n131), .Z(n180) );
  GTECH_NOT U214 ( .A(n124), .Z(n131) );
  GTECH_NAND2 U215 ( .A(n183), .B(n123), .Z(n124) );
  GTECH_NOT U216 ( .A(reset), .Z(n123) );
  GTECH_NOT U217 ( .A(n130), .Z(n189) );
  GTECH_NAND5 U218 ( .A(n127), .B(n190), .C(n183), .D(n104), .E(n118), .Z(n130) );
  GTECH_NOT U219 ( .A(n142), .Z(n183) );
  GTECH_NAND5 U220 ( .A(n136), .B(n141), .C(n143), .D(n107), .E(n105), .Z(n142) );
  GTECH_NOT U221 ( .A(n154), .Z(n143) );
  GTECH_NAND5 U222 ( .A(n191), .B(n151), .C(n152), .D(n110), .E(n109), .Z(n154) );
  GTECH_NOT U223 ( .A(n165), .Z(n152) );
  GTECH_NAND5 U224 ( .A(n192), .B(n193), .C(n163), .D(ss[6]), .E(ss[4]), .Z(
        n165) );
  GTECH_NOT U225 ( .A(n175), .Z(n163) );
  GTECH_NAND5 U226 ( .A(n194), .B(n195), .C(ena), .D(ss[3]), .E(ss[0]), .Z(
        n175) );
  GTECH_NOT U227 ( .A(ss[2]), .Z(n195) );
  GTECH_NOT U228 ( .A(ss[1]), .Z(n194) );
  GTECH_NOT U229 ( .A(ss[7]), .Z(n193) );
  GTECH_NOT U230 ( .A(ss[5]), .Z(n192) );
  GTECH_NOT U231 ( .A(n3), .Z(n151) );
  GTECH_NOT U232 ( .A(n108), .Z(n191) );
  GTECH_NOT U233 ( .A(n4), .Z(n141) );
  GTECH_NOT U234 ( .A(n106), .Z(n136) );
  GTECH_NOT U235 ( .A(n8), .Z(n190) );
  GTECH_NOT U236 ( .A(n103), .Z(n127) );
endmodule

