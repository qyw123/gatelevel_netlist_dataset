
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n127, n129, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n129), .K(n129), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n266) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n129), .K(n129), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n129), .K(n129), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n129), .K(n129), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n129), .K(n129), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n129), .K(n129), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]) );
  GTECH_FJK1S A_reg_15_ ( .J(n129), .K(n129), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n282) );
  GTECH_FJK1S A_reg_14_ ( .J(n129), .K(n129), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n281) );
  GTECH_FJK1S A_reg_13_ ( .J(n129), .K(n129), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n280) );
  GTECH_FJK1S A_reg_12_ ( .J(n129), .K(n129), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n279) );
  GTECH_FJK1S A_reg_11_ ( .J(n129), .K(n129), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n278) );
  GTECH_FJK1S A_reg_10_ ( .J(n129), .K(n129), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n277) );
  GTECH_FJK1S A_reg_9_ ( .J(n129), .K(n129), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n276) );
  GTECH_FJK1S A_reg_8_ ( .J(n129), .K(n129), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n275) );
  GTECH_FJK1S A_reg_7_ ( .J(n129), .K(n129), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n274) );
  GTECH_FJK1S A_reg_6_ ( .J(n129), .K(n129), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n273) );
  GTECH_FJK1S A_reg_5_ ( .J(n129), .K(n129), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n272) );
  GTECH_FJK1S A_reg_4_ ( .J(n129), .K(n129), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n271) );
  GTECH_FJK1S A_reg_3_ ( .J(n129), .K(n129), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n270) );
  GTECH_FJK1S A_reg_2_ ( .J(n129), .K(n129), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n269) );
  GTECH_FJK1S A_reg_1_ ( .J(n129), .K(n129), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n268) );
  GTECH_FJK1S A_reg_0_ ( .J(n129), .K(n129), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n267) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n129), .K(n129), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n129), .K(n129), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n129), .K(n129), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n129), .K(n129), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n129), .K(n129), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n129), .K(n129), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n129), .K(n129), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n129), .K(n129), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n129), .K(n129), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n129), .K(n129), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n129), .K(n129), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n129), .K(n129), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n129), .K(n129), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n129), .K(n129), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n129), .K(n129), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n129), .K(n129), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n129), .K(n129), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n129), .K(n129), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n129), .K(n129), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n129), .K(n129), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n129), .K(n129), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n129), .K(n129), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n129), .K(n129), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n129), .K(n129), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n129), .K(n129), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n129), .K(n129), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n129), .K(n129), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n129), .K(n129), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n129), .K(n129), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n129), .K(n129), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n129), .K(n129), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n129), .K(n129), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n129), .K(n129), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n129), .K(n129), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n129), .K(n129), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n129), .K(n129), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n129), .K(n129), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n129), .K(n129), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n129), .K(n129), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n129), .K(n129), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n129), .K(n129), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n129), .K(n129), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n129), .K(n129), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n129), .K(n129), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n129), .K(n129), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n129), .K(n129), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n129), .K(n129), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n129), .K(n129), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n129), .K(n129), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n129), .K(n129), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n129), .K(n129), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n129), .K(n129), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n129), .K(n129), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n129), .K(n129), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n129), .K(n129), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n129), .K(n129), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n129), .K(n129), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n129), .K(n129), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n129), .K(n129), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n129), .K(n129), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n129), .K(n129), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n129), .K(n129), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n129), .K(n129), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n129), .K(n129), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n129), .K(n129), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n129), .K(n129), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD2 Valid_reg ( .D(N155), .CP(clk), .CD(n127), .Q(Valid) );
  GTECH_ZERO U268 ( .Z(n129) );
  GTECH_ONE U269 ( .Z(n127) );
  GTECH_NOT U270 ( .A(n284), .Z(N99) );
  GTECH_AOI222 U271 ( .A(n285), .B(n286), .C(n287), .D(n288), .E(n289), .F(
        n290), .Z(n284) );
  GTECH_NOT U272 ( .A(n291), .Z(N98) );
  GTECH_AOI222 U273 ( .A(n287), .B(n292), .C(n293), .D(n294), .E(R[15]), .F(
        n295), .Z(n291) );
  GTECH_NAND2 U274 ( .A(n296), .B(n297), .Z(n293) );
  GTECH_AO22 U275 ( .A(n298), .B(n299), .C(R[14]), .D(n295), .Z(N97) );
  GTECH_AO22 U276 ( .A(n298), .B(n300), .C(R[13]), .D(n295), .Z(N96) );
  GTECH_AO22 U277 ( .A(n298), .B(n301), .C(R[12]), .D(n295), .Z(N95) );
  GTECH_AO22 U278 ( .A(n298), .B(n302), .C(R[11]), .D(n295), .Z(N94) );
  GTECH_AO22 U279 ( .A(n298), .B(n303), .C(R[10]), .D(n295), .Z(N93) );
  GTECH_AO22 U280 ( .A(n298), .B(n304), .C(R[9]), .D(n295), .Z(N92) );
  GTECH_AO22 U281 ( .A(n298), .B(n305), .C(R[8]), .D(n295), .Z(N91) );
  GTECH_AO22 U282 ( .A(n298), .B(n306), .C(R[7]), .D(n295), .Z(N90) );
  GTECH_AO22 U283 ( .A(n298), .B(n307), .C(R[6]), .D(n295), .Z(N89) );
  GTECH_AO22 U284 ( .A(n298), .B(n308), .C(R[5]), .D(n295), .Z(N88) );
  GTECH_AO22 U285 ( .A(n298), .B(n309), .C(R[4]), .D(n295), .Z(N87) );
  GTECH_AO22 U286 ( .A(n298), .B(n310), .C(R[3]), .D(n295), .Z(N86) );
  GTECH_AO22 U287 ( .A(n298), .B(n311), .C(R[2]), .D(n295), .Z(N85) );
  GTECH_AO22 U288 ( .A(n298), .B(n312), .C(R[1]), .D(n295), .Z(N84) );
  GTECH_AO22 U289 ( .A(n298), .B(n313), .C(R[0]), .D(n295), .Z(N83) );
  GTECH_AND2 U290 ( .A(M[15]), .B(n295), .Z(N42) );
  GTECH_AND2 U291 ( .A(M[14]), .B(n295), .Z(N39) );
  GTECH_AND2 U292 ( .A(M[13]), .B(n295), .Z(N38) );
  GTECH_AND2 U293 ( .A(M[12]), .B(n295), .Z(N37) );
  GTECH_AND2 U294 ( .A(M[11]), .B(n295), .Z(N36) );
  GTECH_AND2 U295 ( .A(M[10]), .B(n295), .Z(N35) );
  GTECH_AND2 U296 ( .A(M[9]), .B(n295), .Z(N34) );
  GTECH_AND2 U297 ( .A(M[8]), .B(n295), .Z(N33) );
  GTECH_AND2 U298 ( .A(M[7]), .B(n295), .Z(N32) );
  GTECH_AND2 U299 ( .A(M[6]), .B(n295), .Z(N31) );
  GTECH_AND2 U300 ( .A(M[5]), .B(n295), .Z(N30) );
  GTECH_AND2 U301 ( .A(M[4]), .B(n295), .Z(N29) );
  GTECH_AND2 U302 ( .A(M[3]), .B(n295), .Z(N28) );
  GTECH_AND2 U303 ( .A(M[2]), .B(n295), .Z(N27) );
  GTECH_AND2 U304 ( .A(M[1]), .B(n295), .Z(N26) );
  GTECH_AND2 U305 ( .A(M[0]), .B(n295), .Z(N25) );
  GTECH_NOT U306 ( .A(n314), .Z(n295) );
  GTECH_NAND2 U307 ( .A(n314), .B(n315), .Z(N19) );
  GTECH_NAND3 U308 ( .A(n316), .B(n317), .C(n298), .Z(n315) );
  GTECH_NAND3 U309 ( .A(n318), .B(n319), .C(n320), .Z(N18) );
  GTECH_AND2 U310 ( .A(n298), .B(n321), .Z(N17) );
  GTECH_OAI21 U311 ( .A(n8), .B(n322), .C(n316), .Z(n321) );
  GTECH_AND2 U312 ( .A(n298), .B(n323), .Z(N16) );
  GTECH_OAI21 U313 ( .A(n7), .B(n324), .C(n325), .Z(n323) );
  GTECH_NOT U314 ( .A(n326), .Z(N152) );
  GTECH_AOI222 U315 ( .A(n327), .B(n328), .C(n329), .D(n330), .E(n331), .F(
        n332), .Z(n326) );
  GTECH_NAND2 U316 ( .A(n319), .B(n333), .Z(N151) );
  GTECH_NOT U317 ( .A(n334), .Z(N150) );
  GTECH_AOI222 U318 ( .A(n335), .B(n327), .C(n329), .D(n336), .E(n331), .F(
        n337), .Z(n334) );
  GTECH_MUX2 U319 ( .A(n338), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND2 U320 ( .A(n298), .B(n339), .Z(n338) );
  GTECH_NOT U321 ( .A(n340), .Z(N149) );
  GTECH_AOI222 U322 ( .A(n341), .B(n327), .C(n329), .D(n342), .E(n331), .F(
        n343), .Z(n340) );
  GTECH_NOT U323 ( .A(n344), .Z(N148) );
  GTECH_AOI222 U324 ( .A(n345), .B(n327), .C(n329), .D(n346), .E(n331), .F(
        n347), .Z(n344) );
  GTECH_NOT U325 ( .A(n348), .Z(N147) );
  GTECH_AOI222 U326 ( .A(n349), .B(n327), .C(n329), .D(n350), .E(n331), .F(
        n351), .Z(n348) );
  GTECH_NOT U327 ( .A(n352), .Z(N146) );
  GTECH_AOI222 U328 ( .A(n353), .B(n327), .C(n329), .D(n354), .E(n331), .F(
        n355), .Z(n352) );
  GTECH_NOT U329 ( .A(n356), .Z(N145) );
  GTECH_AOI222 U330 ( .A(n357), .B(n327), .C(n329), .D(n358), .E(n331), .F(
        n359), .Z(n356) );
  GTECH_NOT U331 ( .A(n360), .Z(N144) );
  GTECH_AOI222 U332 ( .A(n361), .B(n327), .C(n329), .D(n362), .E(n331), .F(
        n363), .Z(n360) );
  GTECH_NOT U333 ( .A(n364), .Z(N143) );
  GTECH_AOI222 U334 ( .A(n365), .B(n327), .C(n329), .D(n366), .E(n331), .F(
        n367), .Z(n364) );
  GTECH_NOT U335 ( .A(n368), .Z(N142) );
  GTECH_AOI222 U336 ( .A(n369), .B(n327), .C(n329), .D(n370), .E(n331), .F(
        n371), .Z(n368) );
  GTECH_NOT U337 ( .A(n372), .Z(N141) );
  GTECH_AOI222 U338 ( .A(n373), .B(n327), .C(n329), .D(n374), .E(n331), .F(
        n375), .Z(n372) );
  GTECH_NOT U339 ( .A(n376), .Z(N140) );
  GTECH_AOI222 U340 ( .A(n377), .B(n327), .C(n329), .D(n378), .E(n331), .F(
        n379), .Z(n376) );
  GTECH_NOT U341 ( .A(n380), .Z(N14) );
  GTECH_NAND2 U342 ( .A(n298), .B(n266), .Z(n380) );
  GTECH_NOT U343 ( .A(n381), .Z(N139) );
  GTECH_AOI222 U344 ( .A(n382), .B(n327), .C(n329), .D(n383), .E(n331), .F(
        n384), .Z(n381) );
  GTECH_NOT U345 ( .A(n385), .Z(N138) );
  GTECH_AOI222 U346 ( .A(n386), .B(n327), .C(n329), .D(n387), .E(n331), .F(
        n388), .Z(n385) );
  GTECH_NOT U347 ( .A(n389), .Z(N137) );
  GTECH_AOI222 U348 ( .A(n390), .B(n327), .C(n329), .D(n391), .E(n331), .F(
        n392), .Z(n389) );
  GTECH_NOT U349 ( .A(n393), .Z(N136) );
  GTECH_AOI222 U350 ( .A(n327), .B(n286), .C(n329), .D(n288), .E(n331), .F(
        n290), .Z(n393) );
  GTECH_NOT U351 ( .A(n394), .Z(n290) );
  GTECH_XOR2 U352 ( .A(n395), .B(n396), .Z(n394) );
  GTECH_NOT U353 ( .A(n397), .Z(n396) );
  GTECH_NOT U354 ( .A(n398), .Z(n329) );
  GTECH_NOT U355 ( .A(n399), .Z(n286) );
  GTECH_XOR2 U356 ( .A(n395), .B(n400), .Z(n399) );
  GTECH_NOT U357 ( .A(n401), .Z(n400) );
  GTECH_XOR2 U358 ( .A(n288), .B(n268), .Z(n395) );
  GTECH_OAI21 U359 ( .A(n12), .B(n398), .C(n402), .Z(N135) );
  GTECH_OAI21 U360 ( .A(n331), .B(n327), .C(n294), .Z(n402) );
  GTECH_OAI21 U361 ( .A(n12), .B(n403), .C(n397), .Z(n294) );
  GTECH_NOT U362 ( .A(n404), .Z(n327) );
  GTECH_NAND3 U363 ( .A(n28), .B(n405), .C(N155), .Z(n404) );
  GTECH_NOT U364 ( .A(n406), .Z(n331) );
  GTECH_NAND3 U365 ( .A(n10), .B(n407), .C(N155), .Z(n406) );
  GTECH_NAND2 U366 ( .A(n408), .B(N155), .Z(n398) );
  GTECH_XOR2 U367 ( .A(n405), .B(n28), .Z(n408) );
  GTECH_AND2 U368 ( .A(N155), .B(n299), .Z(N134) );
  GTECH_NOT U369 ( .A(n13), .Z(n299) );
  GTECH_AND2 U370 ( .A(N155), .B(n300), .Z(N133) );
  GTECH_NOT U371 ( .A(n14), .Z(n300) );
  GTECH_AND2 U372 ( .A(N155), .B(n301), .Z(N132) );
  GTECH_NOT U373 ( .A(n15), .Z(n301) );
  GTECH_AND2 U374 ( .A(N155), .B(n302), .Z(N131) );
  GTECH_NOT U375 ( .A(n16), .Z(n302) );
  GTECH_AND2 U376 ( .A(N155), .B(n303), .Z(N130) );
  GTECH_NOT U377 ( .A(n17), .Z(n303) );
  GTECH_AND2 U378 ( .A(N155), .B(n304), .Z(N129) );
  GTECH_NOT U379 ( .A(n18), .Z(n304) );
  GTECH_AND2 U380 ( .A(N155), .B(n305), .Z(N128) );
  GTECH_NOT U381 ( .A(n19), .Z(n305) );
  GTECH_AND2 U382 ( .A(N155), .B(n306), .Z(N127) );
  GTECH_NOT U383 ( .A(n20), .Z(n306) );
  GTECH_AND2 U384 ( .A(N155), .B(n307), .Z(N126) );
  GTECH_NOT U385 ( .A(n21), .Z(n307) );
  GTECH_AND2 U386 ( .A(N155), .B(n308), .Z(N125) );
  GTECH_NOT U387 ( .A(n22), .Z(n308) );
  GTECH_AND2 U388 ( .A(N155), .B(n309), .Z(N124) );
  GTECH_NOT U389 ( .A(n23), .Z(n309) );
  GTECH_AND2 U390 ( .A(N155), .B(n310), .Z(N123) );
  GTECH_NOT U391 ( .A(n24), .Z(n310) );
  GTECH_AND2 U392 ( .A(N155), .B(n311), .Z(N122) );
  GTECH_NOT U393 ( .A(n25), .Z(n311) );
  GTECH_AND2 U394 ( .A(N155), .B(n312), .Z(N121) );
  GTECH_NOT U395 ( .A(n26), .Z(n312) );
  GTECH_AND2 U396 ( .A(N155), .B(n313), .Z(N120) );
  GTECH_NOT U397 ( .A(n27), .Z(n313) );
  GTECH_NOT U398 ( .A(n333), .Z(N155) );
  GTECH_NAND4 U399 ( .A(n8), .B(n7), .C(n9), .D(n409), .Z(n333) );
  GTECH_AND3 U400 ( .A(n319), .B(n339), .C(n6), .Z(n409) );
  GTECH_NOT U401 ( .A(n266), .Z(n339) );
  GTECH_NOT U402 ( .A(n410), .Z(N116) );
  GTECH_AOI222 U403 ( .A(n287), .B(n330), .C(n289), .D(n332), .E(n328), .F(
        n285), .Z(n410) );
  GTECH_XOR2 U404 ( .A(n411), .B(n412), .Z(n328) );
  GTECH_ADD_ABC U405 ( .A(n31), .B(n282), .C(n413), .COUT(n412) );
  GTECH_XOR2 U406 ( .A(n414), .B(n411), .Z(n332) );
  GTECH_XOR2 U407 ( .A(A[16]), .B(n30), .Z(n411) );
  GTECH_OAI21 U408 ( .A(n415), .B(n31), .C(n416), .Z(n414) );
  GTECH_OAI21 U409 ( .A(n282), .B(n336), .C(n417), .Z(n416) );
  GTECH_NOT U410 ( .A(n30), .Z(n330) );
  GTECH_NAND2 U411 ( .A(n320), .B(n418), .Z(N115) );
  GTECH_NOT U412 ( .A(N41), .Z(n418) );
  GTECH_NAND2 U413 ( .A(n319), .B(n314), .Z(N41) );
  GTECH_NAND2 U414 ( .A(Ld), .B(n319), .Z(n314) );
  GTECH_NOT U415 ( .A(n419), .Z(N113) );
  GTECH_AOI222 U416 ( .A(n287), .B(n336), .C(n289), .D(n337), .E(n335), .F(
        n285), .Z(n419) );
  GTECH_XOR2 U417 ( .A(n420), .B(n413), .Z(n335) );
  GTECH_ADD_ABC U418 ( .A(n32), .B(n281), .C(n421), .COUT(n413) );
  GTECH_NOT U419 ( .A(n422), .Z(n337) );
  GTECH_XOR2 U420 ( .A(n420), .B(n423), .Z(n422) );
  GTECH_NOT U421 ( .A(n417), .Z(n423) );
  GTECH_OAI21 U422 ( .A(n32), .B(n424), .C(n425), .Z(n417) );
  GTECH_OAI21 U423 ( .A(n281), .B(n342), .C(n426), .Z(n425) );
  GTECH_XOR2 U424 ( .A(n415), .B(n31), .Z(n420) );
  GTECH_NOT U425 ( .A(n282), .Z(n415) );
  GTECH_NOT U426 ( .A(n31), .Z(n336) );
  GTECH_NOT U427 ( .A(n427), .Z(N112) );
  GTECH_AOI222 U428 ( .A(n287), .B(n342), .C(n289), .D(n343), .E(n341), .F(
        n285), .Z(n427) );
  GTECH_XOR2 U429 ( .A(n428), .B(n421), .Z(n341) );
  GTECH_ADD_ABC U430 ( .A(n33), .B(n280), .C(n429), .COUT(n421) );
  GTECH_NOT U431 ( .A(n430), .Z(n343) );
  GTECH_XOR2 U432 ( .A(n428), .B(n431), .Z(n430) );
  GTECH_NOT U433 ( .A(n426), .Z(n431) );
  GTECH_OAI21 U434 ( .A(n33), .B(n432), .C(n433), .Z(n426) );
  GTECH_OAI21 U435 ( .A(n280), .B(n346), .C(n434), .Z(n433) );
  GTECH_XOR2 U436 ( .A(n424), .B(n32), .Z(n428) );
  GTECH_NOT U437 ( .A(n281), .Z(n424) );
  GTECH_NOT U438 ( .A(n32), .Z(n342) );
  GTECH_NOT U439 ( .A(n435), .Z(N111) );
  GTECH_AOI222 U440 ( .A(n287), .B(n346), .C(n289), .D(n347), .E(n345), .F(
        n285), .Z(n435) );
  GTECH_XOR2 U441 ( .A(n436), .B(n429), .Z(n345) );
  GTECH_ADD_ABC U442 ( .A(n34), .B(n279), .C(n437), .COUT(n429) );
  GTECH_NOT U443 ( .A(n438), .Z(n347) );
  GTECH_XOR2 U444 ( .A(n436), .B(n439), .Z(n438) );
  GTECH_NOT U445 ( .A(n434), .Z(n439) );
  GTECH_OAI21 U446 ( .A(n34), .B(n440), .C(n441), .Z(n434) );
  GTECH_OAI21 U447 ( .A(n279), .B(n350), .C(n442), .Z(n441) );
  GTECH_XOR2 U448 ( .A(n432), .B(n33), .Z(n436) );
  GTECH_NOT U449 ( .A(n280), .Z(n432) );
  GTECH_NOT U450 ( .A(n33), .Z(n346) );
  GTECH_NOT U451 ( .A(n443), .Z(N110) );
  GTECH_AOI222 U452 ( .A(n287), .B(n350), .C(n289), .D(n351), .E(n349), .F(
        n285), .Z(n443) );
  GTECH_XOR2 U453 ( .A(n444), .B(n437), .Z(n349) );
  GTECH_ADD_ABC U454 ( .A(n35), .B(n278), .C(n445), .COUT(n437) );
  GTECH_NOT U455 ( .A(n446), .Z(n351) );
  GTECH_XOR2 U456 ( .A(n444), .B(n447), .Z(n446) );
  GTECH_NOT U457 ( .A(n442), .Z(n447) );
  GTECH_OAI21 U458 ( .A(n35), .B(n448), .C(n449), .Z(n442) );
  GTECH_OAI21 U459 ( .A(n278), .B(n354), .C(n450), .Z(n449) );
  GTECH_XOR2 U460 ( .A(n440), .B(n34), .Z(n444) );
  GTECH_NOT U461 ( .A(n279), .Z(n440) );
  GTECH_NOT U462 ( .A(n34), .Z(n350) );
  GTECH_NOT U463 ( .A(n451), .Z(N109) );
  GTECH_AOI222 U464 ( .A(n287), .B(n354), .C(n289), .D(n355), .E(n353), .F(
        n285), .Z(n451) );
  GTECH_XOR2 U465 ( .A(n452), .B(n445), .Z(n353) );
  GTECH_ADD_ABC U466 ( .A(n36), .B(n277), .C(n453), .COUT(n445) );
  GTECH_NOT U467 ( .A(n454), .Z(n355) );
  GTECH_XOR2 U468 ( .A(n452), .B(n455), .Z(n454) );
  GTECH_NOT U469 ( .A(n450), .Z(n455) );
  GTECH_OAI21 U470 ( .A(n36), .B(n456), .C(n457), .Z(n450) );
  GTECH_OAI21 U471 ( .A(n277), .B(n358), .C(n458), .Z(n457) );
  GTECH_XOR2 U472 ( .A(n448), .B(n35), .Z(n452) );
  GTECH_NOT U473 ( .A(n278), .Z(n448) );
  GTECH_NOT U474 ( .A(n35), .Z(n354) );
  GTECH_NOT U475 ( .A(n459), .Z(N108) );
  GTECH_AOI222 U476 ( .A(n287), .B(n358), .C(n289), .D(n359), .E(n357), .F(
        n285), .Z(n459) );
  GTECH_XOR2 U477 ( .A(n460), .B(n453), .Z(n357) );
  GTECH_ADD_ABC U478 ( .A(n37), .B(n276), .C(n461), .COUT(n453) );
  GTECH_NOT U479 ( .A(n462), .Z(n359) );
  GTECH_XOR2 U480 ( .A(n460), .B(n463), .Z(n462) );
  GTECH_NOT U481 ( .A(n458), .Z(n463) );
  GTECH_OAI21 U482 ( .A(n37), .B(n464), .C(n465), .Z(n458) );
  GTECH_OAI21 U483 ( .A(n276), .B(n362), .C(n466), .Z(n465) );
  GTECH_XOR2 U484 ( .A(n456), .B(n36), .Z(n460) );
  GTECH_NOT U485 ( .A(n277), .Z(n456) );
  GTECH_NOT U486 ( .A(n36), .Z(n358) );
  GTECH_NOT U487 ( .A(n467), .Z(N107) );
  GTECH_AOI222 U488 ( .A(n287), .B(n362), .C(n289), .D(n363), .E(n361), .F(
        n285), .Z(n467) );
  GTECH_XOR2 U489 ( .A(n468), .B(n461), .Z(n361) );
  GTECH_ADD_ABC U490 ( .A(n38), .B(n275), .C(n469), .COUT(n461) );
  GTECH_NOT U491 ( .A(n470), .Z(n363) );
  GTECH_XOR2 U492 ( .A(n468), .B(n471), .Z(n470) );
  GTECH_NOT U493 ( .A(n466), .Z(n471) );
  GTECH_OAI21 U494 ( .A(n38), .B(n472), .C(n473), .Z(n466) );
  GTECH_OAI21 U495 ( .A(n275), .B(n366), .C(n474), .Z(n473) );
  GTECH_XOR2 U496 ( .A(n464), .B(n37), .Z(n468) );
  GTECH_NOT U497 ( .A(n276), .Z(n464) );
  GTECH_NOT U498 ( .A(n37), .Z(n362) );
  GTECH_NOT U499 ( .A(n475), .Z(N106) );
  GTECH_AOI222 U500 ( .A(n287), .B(n366), .C(n289), .D(n367), .E(n365), .F(
        n285), .Z(n475) );
  GTECH_XOR2 U501 ( .A(n476), .B(n469), .Z(n365) );
  GTECH_ADD_ABC U502 ( .A(n39), .B(n274), .C(n477), .COUT(n469) );
  GTECH_NOT U503 ( .A(n478), .Z(n367) );
  GTECH_XOR2 U504 ( .A(n476), .B(n479), .Z(n478) );
  GTECH_NOT U505 ( .A(n474), .Z(n479) );
  GTECH_OAI21 U506 ( .A(n39), .B(n480), .C(n481), .Z(n474) );
  GTECH_OAI21 U507 ( .A(n274), .B(n370), .C(n482), .Z(n481) );
  GTECH_XOR2 U508 ( .A(n472), .B(n38), .Z(n476) );
  GTECH_NOT U509 ( .A(n275), .Z(n472) );
  GTECH_NOT U510 ( .A(n38), .Z(n366) );
  GTECH_NOT U511 ( .A(n483), .Z(N105) );
  GTECH_AOI222 U512 ( .A(n287), .B(n370), .C(n289), .D(n371), .E(n369), .F(
        n285), .Z(n483) );
  GTECH_XOR2 U513 ( .A(n484), .B(n477), .Z(n369) );
  GTECH_ADD_ABC U514 ( .A(n40), .B(n273), .C(n485), .COUT(n477) );
  GTECH_NOT U515 ( .A(n486), .Z(n371) );
  GTECH_XOR2 U516 ( .A(n484), .B(n487), .Z(n486) );
  GTECH_NOT U517 ( .A(n482), .Z(n487) );
  GTECH_OAI21 U518 ( .A(n40), .B(n488), .C(n489), .Z(n482) );
  GTECH_OAI21 U519 ( .A(n273), .B(n374), .C(n490), .Z(n489) );
  GTECH_XOR2 U520 ( .A(n480), .B(n39), .Z(n484) );
  GTECH_NOT U521 ( .A(n274), .Z(n480) );
  GTECH_NOT U522 ( .A(n39), .Z(n370) );
  GTECH_NOT U523 ( .A(n491), .Z(N104) );
  GTECH_AOI222 U524 ( .A(n287), .B(n374), .C(n289), .D(n375), .E(n373), .F(
        n285), .Z(n491) );
  GTECH_XOR2 U525 ( .A(n492), .B(n485), .Z(n373) );
  GTECH_ADD_ABC U526 ( .A(n41), .B(n272), .C(n493), .COUT(n485) );
  GTECH_NOT U527 ( .A(n494), .Z(n375) );
  GTECH_XOR2 U528 ( .A(n492), .B(n495), .Z(n494) );
  GTECH_NOT U529 ( .A(n490), .Z(n495) );
  GTECH_OAI21 U530 ( .A(n41), .B(n496), .C(n497), .Z(n490) );
  GTECH_OAI21 U531 ( .A(n272), .B(n378), .C(n498), .Z(n497) );
  GTECH_XOR2 U532 ( .A(n488), .B(n40), .Z(n492) );
  GTECH_NOT U533 ( .A(n273), .Z(n488) );
  GTECH_NOT U534 ( .A(n40), .Z(n374) );
  GTECH_NOT U535 ( .A(n499), .Z(N103) );
  GTECH_AOI222 U536 ( .A(n287), .B(n378), .C(n289), .D(n379), .E(n377), .F(
        n285), .Z(n499) );
  GTECH_XOR2 U537 ( .A(n500), .B(n493), .Z(n377) );
  GTECH_ADD_ABC U538 ( .A(n42), .B(n271), .C(n501), .COUT(n493) );
  GTECH_NOT U539 ( .A(n502), .Z(n379) );
  GTECH_XOR2 U540 ( .A(n500), .B(n503), .Z(n502) );
  GTECH_NOT U541 ( .A(n498), .Z(n503) );
  GTECH_OAI21 U542 ( .A(n42), .B(n504), .C(n505), .Z(n498) );
  GTECH_OAI21 U543 ( .A(n271), .B(n383), .C(n506), .Z(n505) );
  GTECH_XOR2 U544 ( .A(n496), .B(n41), .Z(n500) );
  GTECH_NOT U545 ( .A(n272), .Z(n496) );
  GTECH_NOT U546 ( .A(n41), .Z(n378) );
  GTECH_NOT U547 ( .A(n507), .Z(N102) );
  GTECH_AOI222 U548 ( .A(n287), .B(n383), .C(n289), .D(n384), .E(n382), .F(
        n285), .Z(n507) );
  GTECH_XOR2 U549 ( .A(n508), .B(n501), .Z(n382) );
  GTECH_ADD_ABC U550 ( .A(n43), .B(n270), .C(n509), .COUT(n501) );
  GTECH_NOT U551 ( .A(n510), .Z(n384) );
  GTECH_XOR2 U552 ( .A(n508), .B(n511), .Z(n510) );
  GTECH_NOT U553 ( .A(n506), .Z(n511) );
  GTECH_OAI21 U554 ( .A(n43), .B(n512), .C(n513), .Z(n506) );
  GTECH_OAI21 U555 ( .A(n270), .B(n387), .C(n514), .Z(n513) );
  GTECH_XOR2 U556 ( .A(n504), .B(n42), .Z(n508) );
  GTECH_NOT U557 ( .A(n271), .Z(n504) );
  GTECH_NOT U558 ( .A(n42), .Z(n383) );
  GTECH_NOT U559 ( .A(n515), .Z(N101) );
  GTECH_AOI222 U560 ( .A(n287), .B(n387), .C(n289), .D(n388), .E(n386), .F(
        n285), .Z(n515) );
  GTECH_XOR2 U561 ( .A(n516), .B(n509), .Z(n386) );
  GTECH_ADD_ABC U562 ( .A(n29), .B(n269), .C(n517), .COUT(n509) );
  GTECH_NOT U563 ( .A(n518), .Z(n388) );
  GTECH_XOR2 U564 ( .A(n516), .B(n519), .Z(n518) );
  GTECH_NOT U565 ( .A(n514), .Z(n519) );
  GTECH_OAI21 U566 ( .A(n29), .B(n520), .C(n521), .Z(n514) );
  GTECH_OAI21 U567 ( .A(n269), .B(n391), .C(n522), .Z(n521) );
  GTECH_XOR2 U568 ( .A(n512), .B(n43), .Z(n516) );
  GTECH_NOT U569 ( .A(n270), .Z(n512) );
  GTECH_NOT U570 ( .A(n43), .Z(n387) );
  GTECH_NOT U571 ( .A(n523), .Z(N100) );
  GTECH_AOI222 U572 ( .A(n390), .B(n285), .C(n287), .D(n391), .E(n289), .F(
        n392), .Z(n523) );
  GTECH_NOT U573 ( .A(n524), .Z(n392) );
  GTECH_XOR2 U574 ( .A(n525), .B(n526), .Z(n524) );
  GTECH_NOT U575 ( .A(n522), .Z(n526) );
  GTECH_OAI21 U576 ( .A(n11), .B(n527), .C(n528), .Z(n522) );
  GTECH_OAI21 U577 ( .A(n268), .B(n288), .C(n397), .Z(n528) );
  GTECH_NAND2 U578 ( .A(n12), .B(n403), .Z(n397) );
  GTECH_NOT U579 ( .A(n11), .Z(n288) );
  GTECH_NOT U580 ( .A(n268), .Z(n527) );
  GTECH_NOT U581 ( .A(n297), .Z(n289) );
  GTECH_NAND2 U582 ( .A(N82), .B(n10), .Z(n297) );
  GTECH_NOT U583 ( .A(n529), .Z(N82) );
  GTECH_NOT U584 ( .A(n29), .Z(n391) );
  GTECH_NOT U585 ( .A(n530), .Z(n287) );
  GTECH_MUX2 U586 ( .A(n529), .B(n531), .S(n10), .Z(n530) );
  GTECH_NAND2 U587 ( .A(n28), .B(n298), .Z(n531) );
  GTECH_NAND2 U588 ( .A(n298), .B(n407), .Z(n529) );
  GTECH_NOT U589 ( .A(n28), .Z(n407) );
  GTECH_NOT U590 ( .A(n296), .Z(n285) );
  GTECH_NAND3 U591 ( .A(n298), .B(n405), .C(n28), .Z(n296) );
  GTECH_NOT U592 ( .A(n10), .Z(n405) );
  GTECH_NOT U593 ( .A(n320), .Z(n298) );
  GTECH_OAI21 U594 ( .A(n316), .B(n317), .C(n532), .Z(n320) );
  GTECH_AND2 U595 ( .A(n318), .B(n319), .Z(n532) );
  GTECH_NOT U596 ( .A(Rst), .Z(n319) );
  GTECH_NOT U597 ( .A(Ld), .Z(n318) );
  GTECH_NOT U598 ( .A(n9), .Z(n317) );
  GTECH_NAND2 U599 ( .A(n8), .B(n322), .Z(n316) );
  GTECH_NOT U600 ( .A(n325), .Z(n322) );
  GTECH_NAND2 U601 ( .A(n7), .B(n324), .Z(n325) );
  GTECH_NOT U602 ( .A(n533), .Z(n324) );
  GTECH_NAND2 U603 ( .A(n6), .B(n266), .Z(n533) );
  GTECH_XOR2 U604 ( .A(n525), .B(n517), .Z(n390) );
  GTECH_ADD_ABC U605 ( .A(n268), .B(n11), .C(n401), .COUT(n517) );
  GTECH_NAND2 U606 ( .A(n292), .B(n403), .Z(n401) );
  GTECH_NOT U607 ( .A(n267), .Z(n403) );
  GTECH_NOT U608 ( .A(n12), .Z(n292) );
  GTECH_XOR2 U609 ( .A(n520), .B(n29), .Z(n525) );
  GTECH_NOT U610 ( .A(n269), .Z(n520) );
endmodule

