
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n112, n113, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK2S Cntr_reg_0_ ( .J(n113), .K(n113), .TI(N14), .TE(N18), .CP(clk), 
        .CD(n112), .Q(Cntr[0]), .QN(n337) );
  GTECH_FJK2S Cntr_reg_1_ ( .J(n113), .K(n113), .TI(N15), .TE(N18), .CP(clk), 
        .CD(n112), .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK2S Cntr_reg_2_ ( .J(n113), .K(n113), .TI(N16), .TE(N18), .CP(clk), 
        .CD(n112), .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK2S Cntr_reg_3_ ( .J(n113), .K(n113), .TI(N17), .TE(N18), .CP(clk), 
        .CD(n112), .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK2S Cntr_reg_4_ ( .J(n113), .K(n113), .TI(N19), .TE(N18), .CP(clk), 
        .CD(n112), .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK2S A_reg_16_ ( .J(n113), .K(n113), .TI(N42), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[16]), .QN(n354) );
  GTECH_FJK2S A_reg_15_ ( .J(n113), .K(n113), .TI(N42), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[15]), .QN(n353) );
  GTECH_FJK2S A_reg_14_ ( .J(n113), .K(n113), .TI(N39), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[14]), .QN(n352) );
  GTECH_FJK2S A_reg_13_ ( .J(n113), .K(n113), .TI(N38), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[13]), .QN(n351) );
  GTECH_FJK2S A_reg_12_ ( .J(n113), .K(n113), .TI(N37), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[12]), .QN(n350) );
  GTECH_FJK2S A_reg_11_ ( .J(n113), .K(n113), .TI(N36), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[11]), .QN(n349) );
  GTECH_FJK2S A_reg_10_ ( .J(n113), .K(n113), .TI(N35), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[10]), .QN(n348) );
  GTECH_FJK2S A_reg_9_ ( .J(n113), .K(n113), .TI(N34), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[9]), .QN(n347) );
  GTECH_FJK2S A_reg_8_ ( .J(n113), .K(n113), .TI(N33), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[8]), .QN(n346) );
  GTECH_FJK2S A_reg_7_ ( .J(n113), .K(n113), .TI(N32), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[7]), .QN(n345) );
  GTECH_FJK2S A_reg_6_ ( .J(n113), .K(n113), .TI(N31), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[6]), .QN(n344) );
  GTECH_FJK2S A_reg_5_ ( .J(n113), .K(n113), .TI(N30), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[5]), .QN(n343) );
  GTECH_FJK2S A_reg_4_ ( .J(n113), .K(n113), .TI(N29), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[4]), .QN(n342) );
  GTECH_FJK2S A_reg_3_ ( .J(n113), .K(n113), .TI(N28), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[3]), .QN(n341) );
  GTECH_FJK2S A_reg_2_ ( .J(n113), .K(n113), .TI(N27), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[2]), .QN(n340) );
  GTECH_FJK2S A_reg_1_ ( .J(n113), .K(n113), .TI(N26), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[1]), .QN(n339) );
  GTECH_FJK2S A_reg_0_ ( .J(n113), .K(n113), .TI(N25), .TE(N41), .CP(clk), 
        .CD(n112), .Q(A[0]), .QN(n338) );
  GTECH_FJK2S Prod_reg_0_ ( .J(n113), .K(n113), .TI(N82), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[0]), .QN(n10) );
  GTECH_FJK2S Prod_reg_18_ ( .J(n113), .K(n113), .TI(N100), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK2S Prod_reg_17_ ( .J(n113), .K(n113), .TI(N99), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[17]), .QN(n12) );
  GTECH_FJK2S Prod_reg_16_ ( .J(n113), .K(n113), .TI(N98), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[16]), .QN(n13) );
  GTECH_FJK2S Prod_reg_15_ ( .J(n113), .K(n113), .TI(N97), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[15]), .QN(n14) );
  GTECH_FJK2S Prod_reg_14_ ( .J(n113), .K(n113), .TI(N96), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[14]), .QN(n15) );
  GTECH_FJK2S Prod_reg_13_ ( .J(n113), .K(n113), .TI(N95), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[13]), .QN(n16) );
  GTECH_FJK2S Prod_reg_12_ ( .J(n113), .K(n113), .TI(N94), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[12]), .QN(n17) );
  GTECH_FJK2S Prod_reg_11_ ( .J(n113), .K(n113), .TI(N93), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[11]), .QN(n18) );
  GTECH_FJK2S Prod_reg_10_ ( .J(n113), .K(n113), .TI(N92), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[10]), .QN(n19) );
  GTECH_FJK2S Prod_reg_9_ ( .J(n113), .K(n113), .TI(N91), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[9]), .QN(n20) );
  GTECH_FJK2S Prod_reg_8_ ( .J(n113), .K(n113), .TI(N90), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[8]), .QN(n21) );
  GTECH_FJK2S Prod_reg_7_ ( .J(n113), .K(n113), .TI(N89), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[7]), .QN(n22) );
  GTECH_FJK2S Prod_reg_6_ ( .J(n113), .K(n113), .TI(N88), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[6]), .QN(n23) );
  GTECH_FJK2S Prod_reg_5_ ( .J(n113), .K(n113), .TI(N87), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[5]), .QN(n24) );
  GTECH_FJK2S Prod_reg_4_ ( .J(n113), .K(n113), .TI(N86), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[4]), .QN(n25) );
  GTECH_FJK2S Prod_reg_3_ ( .J(n113), .K(n113), .TI(N85), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[3]), .QN(n26) );
  GTECH_FJK2S Prod_reg_2_ ( .J(n113), .K(n113), .TI(N84), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[2]), .QN(n27) );
  GTECH_FJK2S Prod_reg_1_ ( .J(n113), .K(n113), .TI(N83), .TE(N115), .CP(clk), 
        .CD(n112), .Q(Prod[1]), .QN(n28) );
  GTECH_FJK2S Prod_reg_19_ ( .J(n113), .K(n113), .TI(N101), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK2S Prod_reg_33_ ( .J(n113), .K(n113), .TI(N116), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK2S Prod_reg_32_ ( .J(n113), .K(n113), .TI(N116), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK2S Prod_reg_31_ ( .J(n113), .K(n113), .TI(N113), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK2S Prod_reg_30_ ( .J(n113), .K(n113), .TI(N112), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK2S Prod_reg_29_ ( .J(n113), .K(n113), .TI(N111), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK2S Prod_reg_28_ ( .J(n113), .K(n113), .TI(N110), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK2S Prod_reg_27_ ( .J(n113), .K(n113), .TI(N109), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK2S Prod_reg_26_ ( .J(n113), .K(n113), .TI(N108), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK2S Prod_reg_25_ ( .J(n113), .K(n113), .TI(N107), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK2S Prod_reg_24_ ( .J(n113), .K(n113), .TI(N106), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK2S Prod_reg_23_ ( .J(n113), .K(n113), .TI(N105), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK2S Prod_reg_22_ ( .J(n113), .K(n113), .TI(N104), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK2S Prod_reg_21_ ( .J(n113), .K(n113), .TI(N103), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK2S Prod_reg_20_ ( .J(n113), .K(n113), .TI(N102), .TE(N115), .CP(clk), .CD(n112), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK2S P_reg_31_ ( .J(n113), .K(n113), .TI(N152), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[31]) );
  GTECH_FJK2S P_reg_30_ ( .J(n113), .K(n113), .TI(N150), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[30]) );
  GTECH_FJK2S P_reg_29_ ( .J(n113), .K(n113), .TI(N149), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[29]) );
  GTECH_FJK2S P_reg_28_ ( .J(n113), .K(n113), .TI(N148), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[28]) );
  GTECH_FJK2S P_reg_27_ ( .J(n113), .K(n113), .TI(N147), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[27]) );
  GTECH_FJK2S P_reg_26_ ( .J(n113), .K(n113), .TI(N146), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[26]) );
  GTECH_FJK2S P_reg_25_ ( .J(n113), .K(n113), .TI(N145), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[25]) );
  GTECH_FJK2S P_reg_24_ ( .J(n113), .K(n113), .TI(N144), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[24]) );
  GTECH_FJK2S P_reg_23_ ( .J(n113), .K(n113), .TI(N143), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[23]) );
  GTECH_FJK2S P_reg_22_ ( .J(n113), .K(n113), .TI(N142), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[22]) );
  GTECH_FJK2S P_reg_21_ ( .J(n113), .K(n113), .TI(N141), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[21]) );
  GTECH_FJK2S P_reg_20_ ( .J(n113), .K(n113), .TI(N140), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[20]) );
  GTECH_FJK2S P_reg_19_ ( .J(n113), .K(n113), .TI(N139), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[19]) );
  GTECH_FJK2S P_reg_18_ ( .J(n113), .K(n113), .TI(N138), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[18]) );
  GTECH_FJK2S P_reg_17_ ( .J(n113), .K(n113), .TI(N137), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[17]) );
  GTECH_FJK2S P_reg_16_ ( .J(n113), .K(n113), .TI(N136), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[16]) );
  GTECH_FJK2S P_reg_15_ ( .J(n113), .K(n113), .TI(N135), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[15]) );
  GTECH_FJK2S P_reg_14_ ( .J(n113), .K(n113), .TI(N134), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[14]) );
  GTECH_FJK2S P_reg_13_ ( .J(n113), .K(n113), .TI(N133), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[13]) );
  GTECH_FJK2S P_reg_12_ ( .J(n113), .K(n113), .TI(N132), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[12]) );
  GTECH_FJK2S P_reg_11_ ( .J(n113), .K(n113), .TI(N131), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[11]) );
  GTECH_FJK2S P_reg_10_ ( .J(n113), .K(n113), .TI(N130), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[10]) );
  GTECH_FJK2S P_reg_9_ ( .J(n113), .K(n113), .TI(N129), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[9]) );
  GTECH_FJK2S P_reg_8_ ( .J(n113), .K(n113), .TI(N128), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[8]) );
  GTECH_FJK2S P_reg_7_ ( .J(n113), .K(n113), .TI(N127), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[7]) );
  GTECH_FJK2S P_reg_6_ ( .J(n113), .K(n113), .TI(N126), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[6]) );
  GTECH_FJK2S P_reg_5_ ( .J(n113), .K(n113), .TI(N125), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[5]) );
  GTECH_FJK2S P_reg_4_ ( .J(n113), .K(n113), .TI(N124), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[4]) );
  GTECH_FJK2S P_reg_3_ ( .J(n113), .K(n113), .TI(N123), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[3]) );
  GTECH_FJK2S P_reg_2_ ( .J(n113), .K(n113), .TI(N122), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[2]) );
  GTECH_FJK2S P_reg_1_ ( .J(n113), .K(n113), .TI(N121), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[1]) );
  GTECH_FJK2S P_reg_0_ ( .J(n113), .K(n113), .TI(N120), .TE(N151), .CP(clk), 
        .CD(n112), .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U339 ( .Z(n113) );
  GTECH_ONE U340 ( .Z(n112) );
  GTECH_NOT U341 ( .A(n355), .Z(N99) );
  GTECH_AOI222 U342 ( .A(n356), .B(n357), .C(n358), .D(n359), .E(n360), .F(
        n361), .Z(n355) );
  GTECH_NOT U343 ( .A(n362), .Z(N98) );
  GTECH_AOI222 U344 ( .A(n358), .B(n363), .C(n364), .D(n365), .E(R[15]), .F(
        n366), .Z(n362) );
  GTECH_NAND2 U345 ( .A(n367), .B(n368), .Z(n364) );
  GTECH_OAI2N2 U346 ( .A(n13), .B(n369), .C(R[14]), .D(n366), .Z(N97) );
  GTECH_OAI2N2 U347 ( .A(n14), .B(n369), .C(R[13]), .D(n366), .Z(N96) );
  GTECH_OAI2N2 U348 ( .A(n15), .B(n369), .C(R[12]), .D(n366), .Z(N95) );
  GTECH_OAI2N2 U349 ( .A(n16), .B(n369), .C(R[11]), .D(n366), .Z(N94) );
  GTECH_OAI2N2 U350 ( .A(n17), .B(n369), .C(R[10]), .D(n366), .Z(N93) );
  GTECH_OAI2N2 U351 ( .A(n18), .B(n369), .C(R[9]), .D(n366), .Z(N92) );
  GTECH_OAI2N2 U352 ( .A(n19), .B(n369), .C(R[8]), .D(n366), .Z(N91) );
  GTECH_OAI2N2 U353 ( .A(n20), .B(n369), .C(R[7]), .D(n366), .Z(N90) );
  GTECH_OAI2N2 U354 ( .A(n21), .B(n369), .C(R[6]), .D(n366), .Z(N89) );
  GTECH_OAI2N2 U355 ( .A(n22), .B(n369), .C(R[5]), .D(n366), .Z(N88) );
  GTECH_OAI2N2 U356 ( .A(n23), .B(n369), .C(R[4]), .D(n366), .Z(N87) );
  GTECH_OAI2N2 U357 ( .A(n24), .B(n369), .C(R[3]), .D(n366), .Z(N86) );
  GTECH_OAI2N2 U358 ( .A(n25), .B(n369), .C(R[2]), .D(n366), .Z(N85) );
  GTECH_OAI2N2 U359 ( .A(n26), .B(n369), .C(R[1]), .D(n366), .Z(N84) );
  GTECH_OAI2N2 U360 ( .A(n27), .B(n369), .C(R[0]), .D(n366), .Z(N83) );
  GTECH_AND2 U361 ( .A(M[15]), .B(n366), .Z(N42) );
  GTECH_AND2 U362 ( .A(M[14]), .B(n366), .Z(N39) );
  GTECH_AND2 U363 ( .A(M[13]), .B(n366), .Z(N38) );
  GTECH_AND2 U364 ( .A(M[12]), .B(n366), .Z(N37) );
  GTECH_AND2 U365 ( .A(M[11]), .B(n366), .Z(N36) );
  GTECH_AND2 U366 ( .A(M[10]), .B(n366), .Z(N35) );
  GTECH_AND2 U367 ( .A(M[9]), .B(n366), .Z(N34) );
  GTECH_AND2 U368 ( .A(M[8]), .B(n366), .Z(N33) );
  GTECH_AND2 U369 ( .A(M[7]), .B(n366), .Z(N32) );
  GTECH_AND2 U370 ( .A(M[6]), .B(n366), .Z(N31) );
  GTECH_AND2 U371 ( .A(M[5]), .B(n366), .Z(N30) );
  GTECH_AND2 U372 ( .A(M[4]), .B(n366), .Z(N29) );
  GTECH_AND2 U373 ( .A(M[3]), .B(n366), .Z(N28) );
  GTECH_AND2 U374 ( .A(M[2]), .B(n366), .Z(N27) );
  GTECH_AND2 U375 ( .A(M[1]), .B(n366), .Z(N26) );
  GTECH_AND2 U376 ( .A(M[0]), .B(n366), .Z(N25) );
  GTECH_NOT U377 ( .A(n370), .Z(n366) );
  GTECH_NAND2 U378 ( .A(n370), .B(n371), .Z(N19) );
  GTECH_NAND3 U379 ( .A(n372), .B(n373), .C(n374), .Z(n371) );
  GTECH_NAND3 U380 ( .A(n375), .B(n376), .C(n369), .Z(N18) );
  GTECH_AND2 U381 ( .A(n374), .B(n377), .Z(N17) );
  GTECH_OAI21 U382 ( .A(n8), .B(n378), .C(n372), .Z(n377) );
  GTECH_AND2 U383 ( .A(n374), .B(n379), .Z(N16) );
  GTECH_OAI21 U384 ( .A(n7), .B(n380), .C(n381), .Z(n379) );
  GTECH_NOT U385 ( .A(n382), .Z(N152) );
  GTECH_AOI222 U386 ( .A(n383), .B(n384), .C(n385), .D(n386), .E(n387), .F(
        n388), .Z(n382) );
  GTECH_NAND2 U387 ( .A(n376), .B(n389), .Z(N151) );
  GTECH_NOT U388 ( .A(n390), .Z(N150) );
  GTECH_AOI222 U389 ( .A(n391), .B(n383), .C(n385), .D(n392), .E(n387), .F(
        n393), .Z(n390) );
  GTECH_MUX2 U390 ( .A(n394), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND_NOT U391 ( .A(n374), .B(n337), .Z(n394) );
  GTECH_NOT U392 ( .A(n395), .Z(N149) );
  GTECH_AOI222 U393 ( .A(n396), .B(n383), .C(n385), .D(n397), .E(n387), .F(
        n398), .Z(n395) );
  GTECH_NOT U394 ( .A(n399), .Z(N148) );
  GTECH_AOI222 U395 ( .A(n400), .B(n383), .C(n385), .D(n401), .E(n387), .F(
        n402), .Z(n399) );
  GTECH_NOT U396 ( .A(n403), .Z(N147) );
  GTECH_AOI222 U397 ( .A(n404), .B(n383), .C(n385), .D(n405), .E(n387), .F(
        n406), .Z(n403) );
  GTECH_NOT U398 ( .A(n407), .Z(N146) );
  GTECH_AOI222 U399 ( .A(n408), .B(n383), .C(n385), .D(n409), .E(n387), .F(
        n410), .Z(n407) );
  GTECH_NOT U400 ( .A(n411), .Z(N145) );
  GTECH_AOI222 U401 ( .A(n412), .B(n383), .C(n385), .D(n413), .E(n387), .F(
        n414), .Z(n411) );
  GTECH_NOT U402 ( .A(n415), .Z(N144) );
  GTECH_AOI222 U403 ( .A(n416), .B(n383), .C(n385), .D(n417), .E(n387), .F(
        n418), .Z(n415) );
  GTECH_NOT U404 ( .A(n419), .Z(N143) );
  GTECH_AOI222 U405 ( .A(n420), .B(n383), .C(n385), .D(n421), .E(n387), .F(
        n422), .Z(n419) );
  GTECH_NOT U406 ( .A(n423), .Z(N142) );
  GTECH_AOI222 U407 ( .A(n424), .B(n383), .C(n385), .D(n425), .E(n387), .F(
        n426), .Z(n423) );
  GTECH_NOT U408 ( .A(n427), .Z(N141) );
  GTECH_AOI222 U409 ( .A(n428), .B(n383), .C(n385), .D(n429), .E(n387), .F(
        n430), .Z(n427) );
  GTECH_NOT U410 ( .A(n431), .Z(N140) );
  GTECH_AOI222 U411 ( .A(n432), .B(n383), .C(n385), .D(n433), .E(n387), .F(
        n434), .Z(n431) );
  GTECH_NOT U412 ( .A(n435), .Z(N14) );
  GTECH_NAND2 U413 ( .A(n374), .B(n337), .Z(n435) );
  GTECH_NOT U414 ( .A(n436), .Z(N139) );
  GTECH_AOI222 U415 ( .A(n437), .B(n383), .C(n385), .D(n438), .E(n387), .F(
        n439), .Z(n436) );
  GTECH_NOT U416 ( .A(n440), .Z(N138) );
  GTECH_AOI222 U417 ( .A(n441), .B(n383), .C(n385), .D(n442), .E(n387), .F(
        n443), .Z(n440) );
  GTECH_NOT U418 ( .A(n444), .Z(N137) );
  GTECH_AOI222 U419 ( .A(n445), .B(n383), .C(n385), .D(n446), .E(n387), .F(
        n447), .Z(n444) );
  GTECH_NOT U420 ( .A(n448), .Z(N136) );
  GTECH_AOI222 U421 ( .A(n383), .B(n357), .C(n385), .D(n359), .E(n387), .F(
        n361), .Z(n448) );
  GTECH_NOT U422 ( .A(n449), .Z(n361) );
  GTECH_XOR2 U423 ( .A(n450), .B(n451), .Z(n449) );
  GTECH_NOT U424 ( .A(n452), .Z(n451) );
  GTECH_NOT U425 ( .A(n453), .Z(n385) );
  GTECH_NOT U426 ( .A(n454), .Z(n357) );
  GTECH_XOR2 U427 ( .A(n450), .B(n455), .Z(n454) );
  GTECH_NOT U428 ( .A(n456), .Z(n455) );
  GTECH_XOR2 U429 ( .A(n359), .B(n339), .Z(n450) );
  GTECH_OAI21 U430 ( .A(n12), .B(n453), .C(n457), .Z(N135) );
  GTECH_OAI21 U431 ( .A(n387), .B(n383), .C(n365), .Z(n457) );
  GTECH_OAI21 U432 ( .A(n12), .B(n458), .C(n452), .Z(n365) );
  GTECH_NOT U433 ( .A(n459), .Z(n383) );
  GTECH_NAND3 U434 ( .A(n28), .B(n460), .C(N155), .Z(n459) );
  GTECH_NOT U435 ( .A(n461), .Z(n387) );
  GTECH_NAND3 U436 ( .A(n10), .B(n462), .C(N155), .Z(n461) );
  GTECH_NAND2 U437 ( .A(n463), .B(N155), .Z(n453) );
  GTECH_XOR2 U438 ( .A(n460), .B(n28), .Z(n463) );
  GTECH_AND2 U439 ( .A(N155), .B(n464), .Z(N134) );
  GTECH_NOT U440 ( .A(n13), .Z(n464) );
  GTECH_AND2 U441 ( .A(N155), .B(n465), .Z(N133) );
  GTECH_NOT U442 ( .A(n14), .Z(n465) );
  GTECH_AND2 U443 ( .A(N155), .B(n466), .Z(N132) );
  GTECH_NOT U444 ( .A(n15), .Z(n466) );
  GTECH_AND2 U445 ( .A(N155), .B(n467), .Z(N131) );
  GTECH_NOT U446 ( .A(n16), .Z(n467) );
  GTECH_AND2 U447 ( .A(N155), .B(n468), .Z(N130) );
  GTECH_NOT U448 ( .A(n17), .Z(n468) );
  GTECH_AND2 U449 ( .A(N155), .B(n469), .Z(N129) );
  GTECH_NOT U450 ( .A(n18), .Z(n469) );
  GTECH_AND2 U451 ( .A(N155), .B(n470), .Z(N128) );
  GTECH_NOT U452 ( .A(n19), .Z(n470) );
  GTECH_AND2 U453 ( .A(N155), .B(n471), .Z(N127) );
  GTECH_NOT U454 ( .A(n20), .Z(n471) );
  GTECH_AND2 U455 ( .A(N155), .B(n472), .Z(N126) );
  GTECH_NOT U456 ( .A(n21), .Z(n472) );
  GTECH_AND2 U457 ( .A(N155), .B(n473), .Z(N125) );
  GTECH_NOT U458 ( .A(n22), .Z(n473) );
  GTECH_AND2 U459 ( .A(N155), .B(n474), .Z(N124) );
  GTECH_NOT U460 ( .A(n23), .Z(n474) );
  GTECH_AND2 U461 ( .A(N155), .B(n475), .Z(N123) );
  GTECH_NOT U462 ( .A(n24), .Z(n475) );
  GTECH_AND2 U463 ( .A(N155), .B(n476), .Z(N122) );
  GTECH_NOT U464 ( .A(n25), .Z(n476) );
  GTECH_AND2 U465 ( .A(N155), .B(n477), .Z(N121) );
  GTECH_NOT U466 ( .A(n26), .Z(n477) );
  GTECH_AND2 U467 ( .A(N155), .B(n478), .Z(N120) );
  GTECH_NOT U468 ( .A(n27), .Z(n478) );
  GTECH_NOT U469 ( .A(n389), .Z(N155) );
  GTECH_NAND5 U470 ( .A(n479), .B(n6), .C(n9), .D(n8), .E(n7), .Z(n389) );
  GTECH_NOR2 U471 ( .A(n337), .B(Rst), .Z(n479) );
  GTECH_NOT U472 ( .A(n480), .Z(N116) );
  GTECH_AOI222 U473 ( .A(n358), .B(n386), .C(n360), .D(n388), .E(n384), .F(
        n356), .Z(n480) );
  GTECH_XOR2 U474 ( .A(n481), .B(n482), .Z(n384) );
  GTECH_ADD_ABC U475 ( .A(n353), .B(n31), .C(n483), .COUT(n482) );
  GTECH_XOR2 U476 ( .A(n484), .B(n481), .Z(n388) );
  GTECH_XOR2 U477 ( .A(n386), .B(n354), .Z(n481) );
  GTECH_NAND2 U478 ( .A(n485), .B(n486), .Z(n484) );
  GTECH_OAI21 U479 ( .A(n353), .B(n392), .C(n487), .Z(n486) );
  GTECH_OR_NOT U480 ( .A(n31), .B(n353), .Z(n485) );
  GTECH_NOT U481 ( .A(n30), .Z(n386) );
  GTECH_NAND2 U482 ( .A(n369), .B(n488), .Z(N115) );
  GTECH_NOT U483 ( .A(N41), .Z(n488) );
  GTECH_NAND2 U484 ( .A(n376), .B(n370), .Z(N41) );
  GTECH_NAND2 U485 ( .A(Ld), .B(n376), .Z(n370) );
  GTECH_NOT U486 ( .A(n489), .Z(N113) );
  GTECH_AOI222 U487 ( .A(n358), .B(n392), .C(n360), .D(n393), .E(n391), .F(
        n356), .Z(n489) );
  GTECH_XOR2 U488 ( .A(n490), .B(n483), .Z(n391) );
  GTECH_ADD_ABC U489 ( .A(n352), .B(n32), .C(n491), .COUT(n483) );
  GTECH_NOT U490 ( .A(n492), .Z(n393) );
  GTECH_XOR2 U491 ( .A(n490), .B(n493), .Z(n492) );
  GTECH_NOT U492 ( .A(n487), .Z(n493) );
  GTECH_OAI21 U493 ( .A(n32), .B(n494), .C(n495), .Z(n487) );
  GTECH_OAI21 U494 ( .A(n352), .B(n397), .C(n496), .Z(n495) );
  GTECH_NOT U495 ( .A(n352), .Z(n494) );
  GTECH_XOR2 U496 ( .A(n392), .B(n353), .Z(n490) );
  GTECH_NOT U497 ( .A(n31), .Z(n392) );
  GTECH_NOT U498 ( .A(n497), .Z(N112) );
  GTECH_AOI222 U499 ( .A(n358), .B(n397), .C(n360), .D(n398), .E(n396), .F(
        n356), .Z(n497) );
  GTECH_XOR2 U500 ( .A(n498), .B(n491), .Z(n396) );
  GTECH_ADD_ABC U501 ( .A(n33), .B(n351), .C(n499), .COUT(n491) );
  GTECH_NOT U502 ( .A(n500), .Z(n398) );
  GTECH_XOR2 U503 ( .A(n498), .B(n501), .Z(n500) );
  GTECH_NOT U504 ( .A(n496), .Z(n501) );
  GTECH_OAI21 U505 ( .A(n33), .B(n502), .C(n503), .Z(n496) );
  GTECH_OAI21 U506 ( .A(n351), .B(n401), .C(n504), .Z(n503) );
  GTECH_XOR2 U507 ( .A(n397), .B(n352), .Z(n498) );
  GTECH_NOT U508 ( .A(n32), .Z(n397) );
  GTECH_NOT U509 ( .A(n505), .Z(N111) );
  GTECH_AOI222 U510 ( .A(n358), .B(n401), .C(n360), .D(n402), .E(n400), .F(
        n356), .Z(n505) );
  GTECH_XOR2 U511 ( .A(n506), .B(n499), .Z(n400) );
  GTECH_ADD_ABC U512 ( .A(n34), .B(n350), .C(n507), .COUT(n499) );
  GTECH_NOT U513 ( .A(n508), .Z(n402) );
  GTECH_XOR2 U514 ( .A(n506), .B(n509), .Z(n508) );
  GTECH_NOT U515 ( .A(n504), .Z(n509) );
  GTECH_OAI21 U516 ( .A(n34), .B(n510), .C(n511), .Z(n504) );
  GTECH_OAI21 U517 ( .A(n350), .B(n405), .C(n512), .Z(n511) );
  GTECH_XOR2 U518 ( .A(n502), .B(n33), .Z(n506) );
  GTECH_NOT U519 ( .A(n351), .Z(n502) );
  GTECH_NOT U520 ( .A(n33), .Z(n401) );
  GTECH_NOT U521 ( .A(n513), .Z(N110) );
  GTECH_AOI222 U522 ( .A(n358), .B(n405), .C(n360), .D(n406), .E(n404), .F(
        n356), .Z(n513) );
  GTECH_XOR2 U523 ( .A(n514), .B(n507), .Z(n404) );
  GTECH_ADD_ABC U524 ( .A(n35), .B(n349), .C(n515), .COUT(n507) );
  GTECH_NOT U525 ( .A(n516), .Z(n406) );
  GTECH_XOR2 U526 ( .A(n514), .B(n517), .Z(n516) );
  GTECH_NOT U527 ( .A(n512), .Z(n517) );
  GTECH_OAI21 U528 ( .A(n35), .B(n518), .C(n519), .Z(n512) );
  GTECH_OAI21 U529 ( .A(n349), .B(n409), .C(n520), .Z(n519) );
  GTECH_XOR2 U530 ( .A(n510), .B(n34), .Z(n514) );
  GTECH_NOT U531 ( .A(n350), .Z(n510) );
  GTECH_NOT U532 ( .A(n34), .Z(n405) );
  GTECH_NOT U533 ( .A(n521), .Z(N109) );
  GTECH_AOI222 U534 ( .A(n358), .B(n409), .C(n360), .D(n410), .E(n408), .F(
        n356), .Z(n521) );
  GTECH_XOR2 U535 ( .A(n522), .B(n515), .Z(n408) );
  GTECH_ADD_ABC U536 ( .A(n36), .B(n348), .C(n523), .COUT(n515) );
  GTECH_NOT U537 ( .A(n524), .Z(n410) );
  GTECH_XOR2 U538 ( .A(n522), .B(n525), .Z(n524) );
  GTECH_NOT U539 ( .A(n520), .Z(n525) );
  GTECH_OAI21 U540 ( .A(n36), .B(n526), .C(n527), .Z(n520) );
  GTECH_OAI21 U541 ( .A(n348), .B(n413), .C(n528), .Z(n527) );
  GTECH_XOR2 U542 ( .A(n518), .B(n35), .Z(n522) );
  GTECH_NOT U543 ( .A(n349), .Z(n518) );
  GTECH_NOT U544 ( .A(n35), .Z(n409) );
  GTECH_NOT U545 ( .A(n529), .Z(N108) );
  GTECH_AOI222 U546 ( .A(n358), .B(n413), .C(n360), .D(n414), .E(n412), .F(
        n356), .Z(n529) );
  GTECH_XOR2 U547 ( .A(n530), .B(n523), .Z(n412) );
  GTECH_ADD_ABC U548 ( .A(n37), .B(n347), .C(n531), .COUT(n523) );
  GTECH_NOT U549 ( .A(n532), .Z(n414) );
  GTECH_XOR2 U550 ( .A(n530), .B(n533), .Z(n532) );
  GTECH_NOT U551 ( .A(n528), .Z(n533) );
  GTECH_OAI21 U552 ( .A(n37), .B(n534), .C(n535), .Z(n528) );
  GTECH_OAI21 U553 ( .A(n347), .B(n417), .C(n536), .Z(n535) );
  GTECH_XOR2 U554 ( .A(n526), .B(n36), .Z(n530) );
  GTECH_NOT U555 ( .A(n348), .Z(n526) );
  GTECH_NOT U556 ( .A(n36), .Z(n413) );
  GTECH_NOT U557 ( .A(n537), .Z(N107) );
  GTECH_AOI222 U558 ( .A(n358), .B(n417), .C(n360), .D(n418), .E(n416), .F(
        n356), .Z(n537) );
  GTECH_XOR2 U559 ( .A(n538), .B(n531), .Z(n416) );
  GTECH_ADD_ABC U560 ( .A(n38), .B(n346), .C(n539), .COUT(n531) );
  GTECH_NOT U561 ( .A(n540), .Z(n418) );
  GTECH_XOR2 U562 ( .A(n538), .B(n541), .Z(n540) );
  GTECH_NOT U563 ( .A(n536), .Z(n541) );
  GTECH_OAI21 U564 ( .A(n38), .B(n542), .C(n543), .Z(n536) );
  GTECH_OAI21 U565 ( .A(n346), .B(n421), .C(n544), .Z(n543) );
  GTECH_XOR2 U566 ( .A(n534), .B(n37), .Z(n538) );
  GTECH_NOT U567 ( .A(n347), .Z(n534) );
  GTECH_NOT U568 ( .A(n37), .Z(n417) );
  GTECH_NOT U569 ( .A(n545), .Z(N106) );
  GTECH_AOI222 U570 ( .A(n358), .B(n421), .C(n360), .D(n422), .E(n420), .F(
        n356), .Z(n545) );
  GTECH_XOR2 U571 ( .A(n546), .B(n539), .Z(n420) );
  GTECH_ADD_ABC U572 ( .A(n39), .B(n345), .C(n547), .COUT(n539) );
  GTECH_NOT U573 ( .A(n548), .Z(n422) );
  GTECH_XOR2 U574 ( .A(n546), .B(n549), .Z(n548) );
  GTECH_NOT U575 ( .A(n544), .Z(n549) );
  GTECH_OAI21 U576 ( .A(n39), .B(n550), .C(n551), .Z(n544) );
  GTECH_OAI21 U577 ( .A(n345), .B(n425), .C(n552), .Z(n551) );
  GTECH_XOR2 U578 ( .A(n542), .B(n38), .Z(n546) );
  GTECH_NOT U579 ( .A(n346), .Z(n542) );
  GTECH_NOT U580 ( .A(n38), .Z(n421) );
  GTECH_NOT U581 ( .A(n553), .Z(N105) );
  GTECH_AOI222 U582 ( .A(n358), .B(n425), .C(n360), .D(n426), .E(n424), .F(
        n356), .Z(n553) );
  GTECH_XOR2 U583 ( .A(n554), .B(n547), .Z(n424) );
  GTECH_ADD_ABC U584 ( .A(n40), .B(n344), .C(n555), .COUT(n547) );
  GTECH_NOT U585 ( .A(n556), .Z(n426) );
  GTECH_XOR2 U586 ( .A(n554), .B(n557), .Z(n556) );
  GTECH_NOT U587 ( .A(n552), .Z(n557) );
  GTECH_OAI21 U588 ( .A(n40), .B(n558), .C(n559), .Z(n552) );
  GTECH_OAI21 U589 ( .A(n344), .B(n429), .C(n560), .Z(n559) );
  GTECH_XOR2 U590 ( .A(n550), .B(n39), .Z(n554) );
  GTECH_NOT U591 ( .A(n345), .Z(n550) );
  GTECH_NOT U592 ( .A(n39), .Z(n425) );
  GTECH_NOT U593 ( .A(n561), .Z(N104) );
  GTECH_AOI222 U594 ( .A(n358), .B(n429), .C(n360), .D(n430), .E(n428), .F(
        n356), .Z(n561) );
  GTECH_XOR2 U595 ( .A(n562), .B(n555), .Z(n428) );
  GTECH_ADD_ABC U596 ( .A(n41), .B(n343), .C(n563), .COUT(n555) );
  GTECH_NOT U597 ( .A(n564), .Z(n430) );
  GTECH_XOR2 U598 ( .A(n562), .B(n565), .Z(n564) );
  GTECH_NOT U599 ( .A(n560), .Z(n565) );
  GTECH_OAI21 U600 ( .A(n41), .B(n566), .C(n567), .Z(n560) );
  GTECH_OAI21 U601 ( .A(n343), .B(n433), .C(n568), .Z(n567) );
  GTECH_XOR2 U602 ( .A(n558), .B(n40), .Z(n562) );
  GTECH_NOT U603 ( .A(n344), .Z(n558) );
  GTECH_NOT U604 ( .A(n40), .Z(n429) );
  GTECH_NOT U605 ( .A(n569), .Z(N103) );
  GTECH_AOI222 U606 ( .A(n358), .B(n433), .C(n360), .D(n434), .E(n432), .F(
        n356), .Z(n569) );
  GTECH_XOR2 U607 ( .A(n570), .B(n563), .Z(n432) );
  GTECH_ADD_ABC U608 ( .A(n42), .B(n342), .C(n571), .COUT(n563) );
  GTECH_NOT U609 ( .A(n572), .Z(n434) );
  GTECH_XOR2 U610 ( .A(n570), .B(n573), .Z(n572) );
  GTECH_NOT U611 ( .A(n568), .Z(n573) );
  GTECH_OAI21 U612 ( .A(n42), .B(n574), .C(n575), .Z(n568) );
  GTECH_OAI21 U613 ( .A(n342), .B(n438), .C(n576), .Z(n575) );
  GTECH_XOR2 U614 ( .A(n566), .B(n41), .Z(n570) );
  GTECH_NOT U615 ( .A(n343), .Z(n566) );
  GTECH_NOT U616 ( .A(n41), .Z(n433) );
  GTECH_NOT U617 ( .A(n577), .Z(N102) );
  GTECH_AOI222 U618 ( .A(n358), .B(n438), .C(n360), .D(n439), .E(n437), .F(
        n356), .Z(n577) );
  GTECH_XOR2 U619 ( .A(n578), .B(n571), .Z(n437) );
  GTECH_ADD_ABC U620 ( .A(n43), .B(n341), .C(n579), .COUT(n571) );
  GTECH_NOT U621 ( .A(n580), .Z(n439) );
  GTECH_XOR2 U622 ( .A(n578), .B(n581), .Z(n580) );
  GTECH_NOT U623 ( .A(n576), .Z(n581) );
  GTECH_OAI21 U624 ( .A(n43), .B(n582), .C(n583), .Z(n576) );
  GTECH_OAI21 U625 ( .A(n341), .B(n442), .C(n584), .Z(n583) );
  GTECH_XOR2 U626 ( .A(n574), .B(n42), .Z(n578) );
  GTECH_NOT U627 ( .A(n342), .Z(n574) );
  GTECH_NOT U628 ( .A(n42), .Z(n438) );
  GTECH_NOT U629 ( .A(n585), .Z(N101) );
  GTECH_AOI222 U630 ( .A(n358), .B(n442), .C(n360), .D(n443), .E(n441), .F(
        n356), .Z(n585) );
  GTECH_XOR2 U631 ( .A(n586), .B(n579), .Z(n441) );
  GTECH_ADD_ABC U632 ( .A(n29), .B(n340), .C(n587), .COUT(n579) );
  GTECH_NOT U633 ( .A(n588), .Z(n443) );
  GTECH_XOR2 U634 ( .A(n586), .B(n589), .Z(n588) );
  GTECH_NOT U635 ( .A(n584), .Z(n589) );
  GTECH_OAI21 U636 ( .A(n29), .B(n590), .C(n591), .Z(n584) );
  GTECH_OAI21 U637 ( .A(n340), .B(n446), .C(n592), .Z(n591) );
  GTECH_XOR2 U638 ( .A(n582), .B(n43), .Z(n586) );
  GTECH_NOT U639 ( .A(n341), .Z(n582) );
  GTECH_NOT U640 ( .A(n43), .Z(n442) );
  GTECH_NOT U641 ( .A(n593), .Z(N100) );
  GTECH_AOI222 U642 ( .A(n445), .B(n356), .C(n358), .D(n446), .E(n360), .F(
        n447), .Z(n593) );
  GTECH_NOT U643 ( .A(n594), .Z(n447) );
  GTECH_XOR2 U644 ( .A(n595), .B(n596), .Z(n594) );
  GTECH_NOT U645 ( .A(n592), .Z(n596) );
  GTECH_OAI21 U646 ( .A(n11), .B(n597), .C(n598), .Z(n592) );
  GTECH_OAI21 U647 ( .A(n339), .B(n359), .C(n452), .Z(n598) );
  GTECH_NAND2 U648 ( .A(n12), .B(n458), .Z(n452) );
  GTECH_NOT U649 ( .A(n11), .Z(n359) );
  GTECH_NOT U650 ( .A(n339), .Z(n597) );
  GTECH_NOT U651 ( .A(n368), .Z(n360) );
  GTECH_NAND2 U652 ( .A(N82), .B(n10), .Z(n368) );
  GTECH_NOT U653 ( .A(n599), .Z(N82) );
  GTECH_NOT U654 ( .A(n29), .Z(n446) );
  GTECH_NOT U655 ( .A(n600), .Z(n358) );
  GTECH_MUX2 U656 ( .A(n599), .B(n601), .S(n10), .Z(n600) );
  GTECH_NAND2 U657 ( .A(n28), .B(n374), .Z(n601) );
  GTECH_NAND2 U658 ( .A(n374), .B(n462), .Z(n599) );
  GTECH_NOT U659 ( .A(n28), .Z(n462) );
  GTECH_NOT U660 ( .A(n367), .Z(n356) );
  GTECH_NAND3 U661 ( .A(n374), .B(n460), .C(n28), .Z(n367) );
  GTECH_NOT U662 ( .A(n10), .Z(n460) );
  GTECH_NOT U663 ( .A(n369), .Z(n374) );
  GTECH_OAI21 U664 ( .A(n372), .B(n373), .C(n602), .Z(n369) );
  GTECH_AND2 U665 ( .A(n375), .B(n376), .Z(n602) );
  GTECH_NOT U666 ( .A(Rst), .Z(n376) );
  GTECH_NOT U667 ( .A(Ld), .Z(n375) );
  GTECH_NOT U668 ( .A(n9), .Z(n373) );
  GTECH_NAND2 U669 ( .A(n8), .B(n378), .Z(n372) );
  GTECH_NOT U670 ( .A(n381), .Z(n378) );
  GTECH_NAND2 U671 ( .A(n7), .B(n380), .Z(n381) );
  GTECH_NOT U672 ( .A(n603), .Z(n380) );
  GTECH_NAND2 U673 ( .A(n6), .B(n337), .Z(n603) );
  GTECH_XOR2 U674 ( .A(n595), .B(n587), .Z(n445) );
  GTECH_ADD_ABC U675 ( .A(n339), .B(n11), .C(n456), .COUT(n587) );
  GTECH_NAND2 U676 ( .A(n363), .B(n458), .Z(n456) );
  GTECH_NOT U677 ( .A(n338), .Z(n458) );
  GTECH_NOT U678 ( .A(n12), .Z(n363) );
  GTECH_XOR2 U679 ( .A(n590), .B(n29), .Z(n595) );
  GTECH_NOT U680 ( .A(n340), .Z(n590) );
endmodule

