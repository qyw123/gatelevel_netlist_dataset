
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375;

  GTECH_MUX2 U131 ( .A(n270), .B(n271), .S(n272), .Z(sum[9]) );
  GTECH_XNOR2 U132 ( .A(n273), .B(n274), .Z(n271) );
  GTECH_XNOR2 U133 ( .A(n274), .B(n275), .Z(n270) );
  GTECH_OAI21 U134 ( .A(b[9]), .B(a[9]), .C(n276), .Z(n274) );
  GTECH_OR_NOT U135 ( .A(n277), .B(n278), .Z(sum[8]) );
  GTECH_OAI21 U136 ( .A(n273), .B(n279), .C(n280), .Z(n278) );
  GTECH_MUX2 U137 ( .A(n281), .B(n282), .S(n283), .Z(sum[7]) );
  GTECH_XOR2 U138 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_XNOR2 U139 ( .A(n286), .B(n284), .Z(n281) );
  GTECH_XOR2 U140 ( .A(n287), .B(b[7]), .Z(n284) );
  GTECH_OA22 U141 ( .A(b[6]), .B(n288), .C(a[6]), .D(n289), .Z(n286) );
  GTECH_AND2 U142 ( .A(a[6]), .B(n289), .Z(n288) );
  GTECH_MUX2 U143 ( .A(n290), .B(n291), .S(n283), .Z(sum[6]) );
  GTECH_XOR2 U144 ( .A(n292), .B(n293), .Z(n291) );
  GTECH_XOR2 U145 ( .A(n292), .B(n289), .Z(n290) );
  GTECH_OR_NOT U146 ( .A(n294), .B(n295), .Z(n289) );
  GTECH_OR3 U147 ( .A(n296), .B(n297), .C(n298), .Z(n295) );
  GTECH_NOT U148 ( .A(n299), .Z(n296) );
  GTECH_XOR2 U149 ( .A(a[6]), .B(b[6]), .Z(n292) );
  GTECH_MUX2 U150 ( .A(n300), .B(n301), .S(n302), .Z(sum[5]) );
  GTECH_AND_NOT U151 ( .A(n299), .B(n294), .Z(n302) );
  GTECH_NAND2 U152 ( .A(n303), .B(n304), .Z(n301) );
  GTECH_AO21 U153 ( .A(b[4]), .B(a[4]), .C(n283), .Z(n304) );
  GTECH_AO22 U154 ( .A(b[4]), .B(a[4]), .C(n303), .D(n283), .Z(n300) );
  GTECH_XNOR2 U155 ( .A(n283), .B(n305), .Z(sum[4]) );
  GTECH_MUX2 U156 ( .A(n306), .B(n307), .S(n308), .Z(sum[3]) );
  GTECH_XNOR2 U157 ( .A(n309), .B(n310), .Z(n307) );
  GTECH_AO21 U158 ( .A(n311), .B(n312), .C(n313), .Z(n309) );
  GTECH_XOR2 U159 ( .A(n314), .B(n310), .Z(n306) );
  GTECH_XOR2 U160 ( .A(a[3]), .B(b[3]), .Z(n310) );
  GTECH_MUX2 U161 ( .A(n315), .B(n316), .S(n308), .Z(sum[2]) );
  GTECH_XOR2 U162 ( .A(n311), .B(n317), .Z(n316) );
  GTECH_NOT U163 ( .A(n318), .Z(n311) );
  GTECH_OAI21 U164 ( .A(n319), .B(n320), .C(n321), .Z(n318) );
  GTECH_XNOR2 U165 ( .A(n317), .B(n322), .Z(n315) );
  GTECH_OAI21 U166 ( .A(a[2]), .B(b[2]), .C(n312), .Z(n317) );
  GTECH_MUX2 U167 ( .A(n323), .B(n324), .S(n325), .Z(sum[1]) );
  GTECH_AND_NOT U168 ( .A(n321), .B(n319), .Z(n325) );
  GTECH_AO21 U169 ( .A(n308), .B(n320), .C(n326), .Z(n324) );
  GTECH_OAI21 U170 ( .A(n326), .B(n308), .C(n320), .Z(n323) );
  GTECH_MUX2 U171 ( .A(n327), .B(n328), .S(n329), .Z(sum[15]) );
  GTECH_XNOR2 U172 ( .A(n330), .B(n331), .Z(n328) );
  GTECH_XNOR2 U173 ( .A(n332), .B(n330), .Z(n327) );
  GTECH_XOR2 U174 ( .A(n333), .B(b[15]), .Z(n330) );
  GTECH_OA22 U175 ( .A(a[14]), .B(n334), .C(b[14]), .D(n335), .Z(n332) );
  GTECH_AND2 U176 ( .A(a[14]), .B(n334), .Z(n335) );
  GTECH_MUX2 U177 ( .A(n336), .B(n337), .S(n329), .Z(sum[14]) );
  GTECH_XNOR2 U178 ( .A(n338), .B(n339), .Z(n337) );
  GTECH_XNOR2 U179 ( .A(n338), .B(n334), .Z(n336) );
  GTECH_OAI2N2 U180 ( .A(n340), .B(n341), .C(a[13]), .D(b[13]), .Z(n334) );
  GTECH_XNOR2 U181 ( .A(a[14]), .B(b[14]), .Z(n338) );
  GTECH_MUX2 U182 ( .A(n342), .B(n343), .S(n329), .Z(sum[13]) );
  GTECH_XNOR2 U183 ( .A(n344), .B(n345), .Z(n343) );
  GTECH_XNOR2 U184 ( .A(n344), .B(n341), .Z(n342) );
  GTECH_NOT U185 ( .A(n346), .Z(n341) );
  GTECH_AOI21 U186 ( .A(a[13]), .B(b[13]), .C(n340), .Z(n344) );
  GTECH_OR_NOT U187 ( .A(n347), .B(n348), .Z(sum[12]) );
  GTECH_OAI21 U188 ( .A(n346), .B(n345), .C(n329), .Z(n348) );
  GTECH_MUX2 U189 ( .A(n349), .B(n350), .S(n272), .Z(sum[11]) );
  GTECH_XNOR2 U190 ( .A(n351), .B(n352), .Z(n350) );
  GTECH_AO21 U191 ( .A(n353), .B(n354), .C(n355), .Z(n351) );
  GTECH_XOR2 U192 ( .A(n356), .B(n352), .Z(n349) );
  GTECH_XOR2 U193 ( .A(a[11]), .B(b[11]), .Z(n352) );
  GTECH_MUX2 U194 ( .A(n357), .B(n358), .S(n272), .Z(sum[10]) );
  GTECH_XOR2 U195 ( .A(n353), .B(n359), .Z(n358) );
  GTECH_AND2 U196 ( .A(n360), .B(n276), .Z(n353) );
  GTECH_OAI21 U197 ( .A(a[9]), .B(b[9]), .C(n273), .Z(n360) );
  GTECH_XOR2 U198 ( .A(n359), .B(n361), .Z(n357) );
  GTECH_OAI21 U199 ( .A(a[10]), .B(b[10]), .C(n354), .Z(n359) );
  GTECH_XOR2 U200 ( .A(cin), .B(n362), .Z(sum[0]) );
  GTECH_AO21 U201 ( .A(n329), .B(n363), .C(n347), .Z(cout) );
  GTECH_NOR3 U202 ( .A(n345), .B(n346), .C(n329), .Z(n347) );
  GTECH_AND2 U203 ( .A(b[12]), .B(a[12]), .Z(n346) );
  GTECH_OAI2N2 U204 ( .A(n364), .B(n333), .C(n365), .D(b[15]), .Z(n363) );
  GTECH_OR_NOT U205 ( .A(n331), .B(n333), .Z(n365) );
  GTECH_NOT U206 ( .A(n364), .Z(n331) );
  GTECH_NOT U207 ( .A(a[15]), .Z(n333) );
  GTECH_AOI21 U208 ( .A(n339), .B(a[14]), .C(n366), .Z(n364) );
  GTECH_NOT U209 ( .A(n367), .Z(n366) );
  GTECH_OAI21 U210 ( .A(a[14]), .B(n339), .C(b[14]), .Z(n367) );
  GTECH_OAI2N2 U211 ( .A(n345), .B(n340), .C(a[13]), .D(b[13]), .Z(n339) );
  GTECH_NOR2 U212 ( .A(a[13]), .B(b[13]), .Z(n340) );
  GTECH_NOR2 U213 ( .A(a[12]), .B(b[12]), .Z(n345) );
  GTECH_AO21 U214 ( .A(n280), .B(n368), .C(n277), .Z(n329) );
  GTECH_NOR3 U215 ( .A(n279), .B(n273), .C(n280), .Z(n277) );
  GTECH_AND2 U216 ( .A(b[8]), .B(a[8]), .Z(n273) );
  GTECH_NOT U217 ( .A(n275), .Z(n279) );
  GTECH_ADD_ABC U218 ( .A(n356), .B(a[11]), .C(b[11]), .COUT(n368) );
  GTECH_AOI21 U219 ( .A(n354), .B(n361), .C(n355), .Z(n356) );
  GTECH_NOR2 U220 ( .A(b[10]), .B(a[10]), .Z(n355) );
  GTECH_AND2 U221 ( .A(n369), .B(n276), .Z(n361) );
  GTECH_NAND2 U222 ( .A(b[9]), .B(a[9]), .Z(n276) );
  GTECH_OAI21 U223 ( .A(b[9]), .B(a[9]), .C(n275), .Z(n369) );
  GTECH_OR2 U224 ( .A(b[8]), .B(a[8]), .Z(n275) );
  GTECH_NAND2 U225 ( .A(a[10]), .B(b[10]), .Z(n354) );
  GTECH_NOT U226 ( .A(n272), .Z(n280) );
  GTECH_MUX2 U227 ( .A(n305), .B(n370), .S(n283), .Z(n272) );
  GTECH_MUX2 U228 ( .A(n371), .B(n362), .S(n308), .Z(n283) );
  GTECH_NOT U229 ( .A(cin), .Z(n308) );
  GTECH_AND_NOT U230 ( .A(n320), .B(n326), .Z(n362) );
  GTECH_NAND2 U231 ( .A(b[0]), .B(a[0]), .Z(n320) );
  GTECH_ADD_ABC U232 ( .A(a[3]), .B(n314), .C(b[3]), .COUT(n371) );
  GTECH_AOI21 U233 ( .A(n312), .B(n372), .C(n313), .Z(n314) );
  GTECH_NOR2 U234 ( .A(b[2]), .B(a[2]), .Z(n313) );
  GTECH_NOT U235 ( .A(n322), .Z(n372) );
  GTECH_OAI21 U236 ( .A(n326), .B(n319), .C(n321), .Z(n322) );
  GTECH_NAND2 U237 ( .A(b[1]), .B(a[1]), .Z(n321) );
  GTECH_NOR2 U238 ( .A(a[1]), .B(b[1]), .Z(n319) );
  GTECH_NOR2 U239 ( .A(a[0]), .B(b[0]), .Z(n326) );
  GTECH_NAND2 U240 ( .A(a[2]), .B(b[2]), .Z(n312) );
  GTECH_AOI2N2 U241 ( .A(n373), .B(b[7]), .C(n285), .D(n287), .Z(n370) );
  GTECH_NAND2 U242 ( .A(n287), .B(n285), .Z(n373) );
  GTECH_AOI21 U243 ( .A(n293), .B(a[6]), .C(n374), .Z(n285) );
  GTECH_NOT U244 ( .A(n375), .Z(n374) );
  GTECH_OAI21 U245 ( .A(a[6]), .B(n293), .C(b[6]), .Z(n375) );
  GTECH_AO21 U246 ( .A(n303), .B(n299), .C(n294), .Z(n293) );
  GTECH_AND2 U247 ( .A(b[5]), .B(a[5]), .Z(n294) );
  GTECH_OR2 U248 ( .A(b[5]), .B(a[5]), .Z(n299) );
  GTECH_OR_NOT U249 ( .A(a[4]), .B(n297), .Z(n303) );
  GTECH_NOT U250 ( .A(b[4]), .Z(n297) );
  GTECH_NOT U251 ( .A(a[7]), .Z(n287) );
  GTECH_XOR2 U252 ( .A(n298), .B(b[4]), .Z(n305) );
  GTECH_NOT U253 ( .A(a[4]), .Z(n298) );
endmodule

