
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376;

  GTECH_MUX2 U140 ( .A(n279), .B(n280), .S(n281), .Z(sum[9]) );
  GTECH_XNOR2 U141 ( .A(n282), .B(n283), .Z(n280) );
  GTECH_XNOR2 U142 ( .A(n284), .B(n283), .Z(n279) );
  GTECH_OAI21 U143 ( .A(a[9]), .B(b[9]), .C(n285), .Z(n283) );
  GTECH_NOT U144 ( .A(n286), .Z(n284) );
  GTECH_AO21 U145 ( .A(n287), .B(n288), .C(n289), .Z(sum[8]) );
  GTECH_OR_NOT U146 ( .A(n286), .B(n290), .Z(n287) );
  GTECH_MUX2 U147 ( .A(n291), .B(n292), .S(n293), .Z(sum[7]) );
  GTECH_XOR2 U148 ( .A(n294), .B(n295), .Z(n292) );
  GTECH_XNOR2 U149 ( .A(n294), .B(n296), .Z(n291) );
  GTECH_AOI21 U150 ( .A(n297), .B(n298), .C(n299), .Z(n296) );
  GTECH_XOR2 U151 ( .A(a[7]), .B(b[7]), .Z(n294) );
  GTECH_MUX2 U152 ( .A(n300), .B(n301), .S(n293), .Z(sum[6]) );
  GTECH_XNOR2 U153 ( .A(n302), .B(n303), .Z(n301) );
  GTECH_XNOR2 U154 ( .A(n302), .B(n297), .Z(n300) );
  GTECH_AO21 U155 ( .A(n304), .B(n305), .C(n306), .Z(n297) );
  GTECH_OR_NOT U156 ( .A(n299), .B(n298), .Z(n302) );
  GTECH_MUX2 U157 ( .A(n307), .B(n308), .S(n309), .Z(sum[5]) );
  GTECH_AND_NOT U158 ( .A(n304), .B(n306), .Z(n309) );
  GTECH_OAI21 U159 ( .A(n305), .B(n293), .C(n310), .Z(n308) );
  GTECH_AO21 U160 ( .A(n310), .B(n293), .C(n305), .Z(n307) );
  GTECH_XNOR2 U161 ( .A(n293), .B(n311), .Z(sum[4]) );
  GTECH_MUX2 U162 ( .A(n312), .B(n313), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U163 ( .A(n314), .B(n315), .Z(n313) );
  GTECH_XOR2 U164 ( .A(n316), .B(n314), .Z(n312) );
  GTECH_XOR2 U165 ( .A(a[3]), .B(b[3]), .Z(n314) );
  GTECH_OA22 U166 ( .A(b[2]), .B(n317), .C(a[2]), .D(n318), .Z(n316) );
  GTECH_AND2 U167 ( .A(n318), .B(a[2]), .Z(n317) );
  GTECH_MUX2 U168 ( .A(n319), .B(n320), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U169 ( .A(n321), .B(n322), .Z(n320) );
  GTECH_XNOR2 U170 ( .A(n321), .B(n318), .Z(n319) );
  GTECH_AO21 U171 ( .A(n323), .B(n324), .C(n325), .Z(n318) );
  GTECH_XNOR2 U172 ( .A(a[2]), .B(b[2]), .Z(n321) );
  GTECH_MUX2 U173 ( .A(n326), .B(n327), .S(n328), .Z(sum[1]) );
  GTECH_AND_NOT U174 ( .A(n323), .B(n325), .Z(n328) );
  GTECH_OAI21 U175 ( .A(cin), .B(n324), .C(n329), .Z(n327) );
  GTECH_AO21 U176 ( .A(n329), .B(cin), .C(n324), .Z(n326) );
  GTECH_MUX2 U177 ( .A(n330), .B(n331), .S(n332), .Z(sum[15]) );
  GTECH_XNOR2 U178 ( .A(n333), .B(n334), .Z(n331) );
  GTECH_XNOR2 U179 ( .A(n335), .B(n333), .Z(n330) );
  GTECH_XNOR2 U180 ( .A(a[15]), .B(b[15]), .Z(n333) );
  GTECH_ADD_ABC U181 ( .A(a[14]), .B(n336), .C(b[14]), .COUT(n335) );
  GTECH_MUX2 U182 ( .A(n337), .B(n338), .S(n332), .Z(sum[14]) );
  GTECH_XOR2 U183 ( .A(n339), .B(n340), .Z(n338) );
  GTECH_XOR2 U184 ( .A(n336), .B(n340), .Z(n337) );
  GTECH_XOR2 U185 ( .A(a[14]), .B(b[14]), .Z(n340) );
  GTECH_AOI21 U186 ( .A(n341), .B(n342), .C(n343), .Z(n336) );
  GTECH_MUX2 U187 ( .A(n344), .B(n345), .S(n332), .Z(sum[13]) );
  GTECH_XOR2 U188 ( .A(n346), .B(n347), .Z(n345) );
  GTECH_XNOR2 U189 ( .A(n348), .B(n347), .Z(n344) );
  GTECH_OAI21 U190 ( .A(a[13]), .B(b[13]), .C(n341), .Z(n347) );
  GTECH_AO21 U191 ( .A(n332), .B(n349), .C(n350), .Z(sum[12]) );
  GTECH_OR_NOT U192 ( .A(n346), .B(n342), .Z(n349) );
  GTECH_NOT U193 ( .A(n348), .Z(n342) );
  GTECH_MUX2 U194 ( .A(n351), .B(n352), .S(n281), .Z(sum[11]) );
  GTECH_XOR2 U195 ( .A(n353), .B(n354), .Z(n352) );
  GTECH_ADD_ABC U196 ( .A(a[10]), .B(n355), .C(b[10]), .COUT(n353) );
  GTECH_XOR2 U197 ( .A(n354), .B(n356), .Z(n351) );
  GTECH_XOR2 U198 ( .A(a[11]), .B(b[11]), .Z(n354) );
  GTECH_MUX2 U199 ( .A(n357), .B(n358), .S(n281), .Z(sum[10]) );
  GTECH_XOR2 U200 ( .A(n355), .B(n359), .Z(n358) );
  GTECH_AOI21 U201 ( .A(n285), .B(n290), .C(n360), .Z(n355) );
  GTECH_NOT U202 ( .A(n282), .Z(n290) );
  GTECH_XOR2 U203 ( .A(n361), .B(n359), .Z(n357) );
  GTECH_XOR2 U204 ( .A(a[10]), .B(b[10]), .Z(n359) );
  GTECH_AO21 U205 ( .A(n362), .B(cin), .C(n363), .Z(sum[0]) );
  GTECH_OR2 U206 ( .A(n324), .B(n364), .Z(n362) );
  GTECH_AO21 U207 ( .A(n332), .B(n365), .C(n350), .Z(cout) );
  GTECH_NOR3 U208 ( .A(n346), .B(n348), .C(n332), .Z(n350) );
  GTECH_AND2 U209 ( .A(b[12]), .B(a[12]), .Z(n348) );
  GTECH_AO22 U210 ( .A(n334), .B(a[15]), .C(n366), .D(b[15]), .Z(n365) );
  GTECH_OR2 U211 ( .A(n334), .B(a[15]), .Z(n366) );
  GTECH_ADD_ABC U212 ( .A(a[14]), .B(n339), .C(b[14]), .COUT(n334) );
  GTECH_AOI21 U213 ( .A(n341), .B(n346), .C(n343), .Z(n339) );
  GTECH_AND_NOT U214 ( .A(n367), .B(b[13]), .Z(n343) );
  GTECH_NOR2 U215 ( .A(a[12]), .B(b[12]), .Z(n346) );
  GTECH_OR_NOT U216 ( .A(n367), .B(b[13]), .Z(n341) );
  GTECH_NOT U217 ( .A(a[13]), .Z(n367) );
  GTECH_AO21 U218 ( .A(n368), .B(n288), .C(n289), .Z(n332) );
  GTECH_NOR3 U219 ( .A(n286), .B(n282), .C(n288), .Z(n289) );
  GTECH_AND2 U220 ( .A(b[8]), .B(a[8]), .Z(n282) );
  GTECH_NOT U221 ( .A(n281), .Z(n288) );
  GTECH_MUX2 U222 ( .A(n311), .B(n369), .S(n293), .Z(n281) );
  GTECH_AO21 U223 ( .A(n370), .B(cin), .C(n363), .Z(n293) );
  GTECH_NOR3 U224 ( .A(n364), .B(cin), .C(n324), .Z(n363) );
  GTECH_AND2 U225 ( .A(a[0]), .B(b[0]), .Z(n324) );
  GTECH_NOT U226 ( .A(n329), .Z(n364) );
  GTECH_AO22 U227 ( .A(n315), .B(a[3]), .C(n371), .D(b[3]), .Z(n370) );
  GTECH_OR2 U228 ( .A(a[3]), .B(n315), .Z(n371) );
  GTECH_AO21 U229 ( .A(n322), .B(a[2]), .C(n372), .Z(n315) );
  GTECH_NOT U230 ( .A(n373), .Z(n372) );
  GTECH_OAI21 U231 ( .A(a[2]), .B(n322), .C(b[2]), .Z(n373) );
  GTECH_AO21 U232 ( .A(n323), .B(n329), .C(n325), .Z(n322) );
  GTECH_AND2 U233 ( .A(b[1]), .B(a[1]), .Z(n325) );
  GTECH_OR2 U234 ( .A(a[0]), .B(b[0]), .Z(n329) );
  GTECH_OR2 U235 ( .A(a[1]), .B(b[1]), .Z(n323) );
  GTECH_AOI22 U236 ( .A(n374), .B(b[7]), .C(n295), .D(a[7]), .Z(n369) );
  GTECH_OR2 U237 ( .A(a[7]), .B(n295), .Z(n374) );
  GTECH_AO21 U238 ( .A(n298), .B(n303), .C(n299), .Z(n295) );
  GTECH_AND2 U239 ( .A(a[6]), .B(b[6]), .Z(n299) );
  GTECH_AO21 U240 ( .A(n310), .B(n304), .C(n306), .Z(n303) );
  GTECH_AND2 U241 ( .A(b[5]), .B(a[5]), .Z(n306) );
  GTECH_OR2 U242 ( .A(a[5]), .B(b[5]), .Z(n304) );
  GTECH_OR2 U243 ( .A(a[6]), .B(b[6]), .Z(n298) );
  GTECH_OR_NOT U244 ( .A(n305), .B(n310), .Z(n311) );
  GTECH_OR2 U245 ( .A(a[4]), .B(b[4]), .Z(n310) );
  GTECH_AND2 U246 ( .A(a[4]), .B(b[4]), .Z(n305) );
  GTECH_AO22 U247 ( .A(n375), .B(b[11]), .C(n356), .D(a[11]), .Z(n368) );
  GTECH_OR2 U248 ( .A(a[11]), .B(n356), .Z(n375) );
  GTECH_ADD_ABC U249 ( .A(n361), .B(a[10]), .C(b[10]), .COUT(n356) );
  GTECH_AOI21 U250 ( .A(n285), .B(n286), .C(n360), .Z(n361) );
  GTECH_AND_NOT U251 ( .A(n376), .B(b[9]), .Z(n360) );
  GTECH_NOR2 U252 ( .A(a[8]), .B(b[8]), .Z(n286) );
  GTECH_OR_NOT U253 ( .A(n376), .B(b[9]), .Z(n285) );
  GTECH_NOT U254 ( .A(a[9]), .Z(n376) );
endmodule

