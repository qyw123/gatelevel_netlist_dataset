
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n112, n114, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n114), .K(n114), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n251) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n114), .K(n114), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n114), .K(n114), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n114), .K(n114), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n114), .K(n114), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n114), .K(n114), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]) );
  GTECH_FJK1S A_reg_15_ ( .J(n114), .K(n114), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n267) );
  GTECH_FJK1S A_reg_14_ ( .J(n114), .K(n114), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n266) );
  GTECH_FJK1S A_reg_13_ ( .J(n114), .K(n114), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n265) );
  GTECH_FJK1S A_reg_12_ ( .J(n114), .K(n114), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n264) );
  GTECH_FJK1S A_reg_11_ ( .J(n114), .K(n114), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n263) );
  GTECH_FJK1S A_reg_10_ ( .J(n114), .K(n114), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n262) );
  GTECH_FJK1S A_reg_9_ ( .J(n114), .K(n114), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n261) );
  GTECH_FJK1S A_reg_8_ ( .J(n114), .K(n114), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n260) );
  GTECH_FJK1S A_reg_7_ ( .J(n114), .K(n114), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n259) );
  GTECH_FJK1S A_reg_6_ ( .J(n114), .K(n114), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n258) );
  GTECH_FJK1S A_reg_5_ ( .J(n114), .K(n114), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n257) );
  GTECH_FJK1S A_reg_4_ ( .J(n114), .K(n114), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n256) );
  GTECH_FJK1S A_reg_3_ ( .J(n114), .K(n114), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n255) );
  GTECH_FJK1S A_reg_2_ ( .J(n114), .K(n114), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n254) );
  GTECH_FJK1S A_reg_1_ ( .J(n114), .K(n114), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n253) );
  GTECH_FJK1S A_reg_0_ ( .J(n114), .K(n114), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n252) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n114), .K(n114), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n114), .K(n114), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n114), .K(n114), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n114), .K(n114), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n114), .K(n114), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n114), .K(n114), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n114), .K(n114), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n114), .K(n114), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n114), .K(n114), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n114), .K(n114), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n114), .K(n114), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n114), .K(n114), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n114), .K(n114), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n114), .K(n114), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n114), .K(n114), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n114), .K(n114), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n114), .K(n114), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n114), .K(n114), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n114), .K(n114), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n114), .K(n114), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n114), .K(n114), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n114), .K(n114), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n114), .K(n114), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n114), .K(n114), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n114), .K(n114), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n114), .K(n114), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n114), .K(n114), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n114), .K(n114), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n114), .K(n114), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n114), .K(n114), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n114), .K(n114), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n114), .K(n114), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n114), .K(n114), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n114), .K(n114), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n114), .K(n114), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n114), .K(n114), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n114), .K(n114), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n114), .K(n114), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n114), .K(n114), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n114), .K(n114), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n114), .K(n114), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n114), .K(n114), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n114), .K(n114), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n114), .K(n114), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n114), .K(n114), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n114), .K(n114), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n114), .K(n114), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n114), .K(n114), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n114), .K(n114), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n114), .K(n114), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n114), .K(n114), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n114), .K(n114), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n114), .K(n114), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n114), .K(n114), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n114), .K(n114), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n114), .K(n114), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n114), .K(n114), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n114), .K(n114), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n114), .K(n114), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n114), .K(n114), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n114), .K(n114), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n114), .K(n114), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n114), .K(n114), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n114), .K(n114), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n114), .K(n114), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n114), .K(n114), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD2 Valid_reg ( .D(N155), .CP(clk), .CD(n112), .Q(Valid) );
  GTECH_ZERO U253 ( .Z(n114) );
  GTECH_ONE U254 ( .Z(n112) );
  GTECH_NOT U255 ( .A(n269), .Z(N99) );
  GTECH_AOI222 U256 ( .A(n270), .B(n271), .C(n272), .D(n273), .E(n274), .F(
        n275), .Z(n269) );
  GTECH_NOT U257 ( .A(n276), .Z(N98) );
  GTECH_AOI222 U258 ( .A(n272), .B(n277), .C(n278), .D(n279), .E(R[15]), .F(
        n280), .Z(n276) );
  GTECH_NAND2 U259 ( .A(n281), .B(n282), .Z(n278) );
  GTECH_OAI2N2 U260 ( .A(n13), .B(n283), .C(R[14]), .D(n280), .Z(N97) );
  GTECH_OAI2N2 U261 ( .A(n14), .B(n283), .C(R[13]), .D(n280), .Z(N96) );
  GTECH_OAI2N2 U262 ( .A(n15), .B(n283), .C(R[12]), .D(n280), .Z(N95) );
  GTECH_OAI2N2 U263 ( .A(n16), .B(n283), .C(R[11]), .D(n280), .Z(N94) );
  GTECH_OAI2N2 U264 ( .A(n17), .B(n283), .C(R[10]), .D(n280), .Z(N93) );
  GTECH_OAI2N2 U265 ( .A(n18), .B(n283), .C(R[9]), .D(n280), .Z(N92) );
  GTECH_OAI2N2 U266 ( .A(n19), .B(n283), .C(R[8]), .D(n280), .Z(N91) );
  GTECH_OAI2N2 U267 ( .A(n20), .B(n283), .C(R[7]), .D(n280), .Z(N90) );
  GTECH_OAI2N2 U268 ( .A(n21), .B(n283), .C(R[6]), .D(n280), .Z(N89) );
  GTECH_OAI2N2 U269 ( .A(n22), .B(n283), .C(R[5]), .D(n280), .Z(N88) );
  GTECH_OAI2N2 U270 ( .A(n23), .B(n283), .C(R[4]), .D(n280), .Z(N87) );
  GTECH_OAI2N2 U271 ( .A(n24), .B(n283), .C(R[3]), .D(n280), .Z(N86) );
  GTECH_OAI2N2 U272 ( .A(n25), .B(n283), .C(R[2]), .D(n280), .Z(N85) );
  GTECH_OAI2N2 U273 ( .A(n26), .B(n283), .C(R[1]), .D(n280), .Z(N84) );
  GTECH_OAI2N2 U274 ( .A(n27), .B(n283), .C(R[0]), .D(n280), .Z(N83) );
  GTECH_AND2 U275 ( .A(M[15]), .B(n280), .Z(N42) );
  GTECH_AND2 U276 ( .A(M[14]), .B(n280), .Z(N39) );
  GTECH_AND2 U277 ( .A(M[13]), .B(n280), .Z(N38) );
  GTECH_AND2 U278 ( .A(M[12]), .B(n280), .Z(N37) );
  GTECH_AND2 U279 ( .A(M[11]), .B(n280), .Z(N36) );
  GTECH_AND2 U280 ( .A(M[10]), .B(n280), .Z(N35) );
  GTECH_AND2 U281 ( .A(M[9]), .B(n280), .Z(N34) );
  GTECH_AND2 U282 ( .A(M[8]), .B(n280), .Z(N33) );
  GTECH_AND2 U283 ( .A(M[7]), .B(n280), .Z(N32) );
  GTECH_AND2 U284 ( .A(M[6]), .B(n280), .Z(N31) );
  GTECH_AND2 U285 ( .A(M[5]), .B(n280), .Z(N30) );
  GTECH_AND2 U286 ( .A(M[4]), .B(n280), .Z(N29) );
  GTECH_AND2 U287 ( .A(M[3]), .B(n280), .Z(N28) );
  GTECH_AND2 U288 ( .A(M[2]), .B(n280), .Z(N27) );
  GTECH_AND2 U289 ( .A(M[1]), .B(n280), .Z(N26) );
  GTECH_AND2 U290 ( .A(M[0]), .B(n280), .Z(N25) );
  GTECH_NOT U291 ( .A(n284), .Z(n280) );
  GTECH_NAND2 U292 ( .A(n284), .B(n285), .Z(N19) );
  GTECH_NAND3 U293 ( .A(n286), .B(n287), .C(n288), .Z(n285) );
  GTECH_NAND3 U294 ( .A(n289), .B(n290), .C(n283), .Z(N18) );
  GTECH_AND2 U295 ( .A(n288), .B(n291), .Z(N17) );
  GTECH_OAI21 U296 ( .A(n8), .B(n292), .C(n286), .Z(n291) );
  GTECH_AND2 U297 ( .A(n288), .B(n293), .Z(N16) );
  GTECH_OAI21 U298 ( .A(n7), .B(n294), .C(n295), .Z(n293) );
  GTECH_NOT U299 ( .A(n296), .Z(N152) );
  GTECH_AOI222 U300 ( .A(n297), .B(n298), .C(n299), .D(n300), .E(n301), .F(
        n302), .Z(n296) );
  GTECH_NAND2 U301 ( .A(n290), .B(n303), .Z(N151) );
  GTECH_NOT U302 ( .A(n304), .Z(N150) );
  GTECH_AOI222 U303 ( .A(n305), .B(n297), .C(n299), .D(n306), .E(n301), .F(
        n307), .Z(n304) );
  GTECH_OAI21 U304 ( .A(n308), .B(n309), .C(n310), .Z(N15) );
  GTECH_NAND3 U305 ( .A(n288), .B(n311), .C(n308), .Z(n310) );
  GTECH_NOT U306 ( .A(n6), .Z(n308) );
  GTECH_NOT U307 ( .A(n312), .Z(N149) );
  GTECH_AOI222 U308 ( .A(n313), .B(n297), .C(n299), .D(n314), .E(n301), .F(
        n315), .Z(n312) );
  GTECH_NOT U309 ( .A(n316), .Z(N148) );
  GTECH_AOI222 U310 ( .A(n317), .B(n297), .C(n299), .D(n318), .E(n301), .F(
        n319), .Z(n316) );
  GTECH_NOT U311 ( .A(n320), .Z(N147) );
  GTECH_AOI222 U312 ( .A(n321), .B(n297), .C(n299), .D(n322), .E(n301), .F(
        n323), .Z(n320) );
  GTECH_NOT U313 ( .A(n324), .Z(N146) );
  GTECH_AOI222 U314 ( .A(n325), .B(n297), .C(n299), .D(n326), .E(n301), .F(
        n327), .Z(n324) );
  GTECH_NOT U315 ( .A(n328), .Z(N145) );
  GTECH_AOI222 U316 ( .A(n329), .B(n297), .C(n299), .D(n330), .E(n301), .F(
        n331), .Z(n328) );
  GTECH_NOT U317 ( .A(n332), .Z(N144) );
  GTECH_AOI222 U318 ( .A(n333), .B(n297), .C(n299), .D(n334), .E(n301), .F(
        n335), .Z(n332) );
  GTECH_NOT U319 ( .A(n336), .Z(N143) );
  GTECH_AOI222 U320 ( .A(n337), .B(n297), .C(n299), .D(n338), .E(n301), .F(
        n339), .Z(n336) );
  GTECH_NOT U321 ( .A(n340), .Z(N142) );
  GTECH_AOI222 U322 ( .A(n341), .B(n297), .C(n299), .D(n342), .E(n301), .F(
        n343), .Z(n340) );
  GTECH_NOT U323 ( .A(n344), .Z(N141) );
  GTECH_AOI222 U324 ( .A(n345), .B(n297), .C(n299), .D(n346), .E(n301), .F(
        n347), .Z(n344) );
  GTECH_NOT U325 ( .A(n348), .Z(N140) );
  GTECH_AOI222 U326 ( .A(n349), .B(n297), .C(n299), .D(n350), .E(n301), .F(
        n351), .Z(n348) );
  GTECH_NOT U327 ( .A(n309), .Z(N14) );
  GTECH_NAND2 U328 ( .A(n288), .B(n251), .Z(n309) );
  GTECH_NOT U329 ( .A(n352), .Z(N139) );
  GTECH_AOI222 U330 ( .A(n353), .B(n297), .C(n299), .D(n354), .E(n301), .F(
        n355), .Z(n352) );
  GTECH_NOT U331 ( .A(n356), .Z(N138) );
  GTECH_AOI222 U332 ( .A(n357), .B(n297), .C(n299), .D(n358), .E(n301), .F(
        n359), .Z(n356) );
  GTECH_NOT U333 ( .A(n360), .Z(N137) );
  GTECH_AOI222 U334 ( .A(n361), .B(n297), .C(n299), .D(n362), .E(n301), .F(
        n363), .Z(n360) );
  GTECH_NOT U335 ( .A(n364), .Z(N136) );
  GTECH_AOI222 U336 ( .A(n297), .B(n271), .C(n299), .D(n273), .E(n301), .F(
        n275), .Z(n364) );
  GTECH_NOT U337 ( .A(n365), .Z(n275) );
  GTECH_XOR2 U338 ( .A(n366), .B(n367), .Z(n365) );
  GTECH_NOT U339 ( .A(n368), .Z(n367) );
  GTECH_NOT U340 ( .A(n369), .Z(n299) );
  GTECH_NOT U341 ( .A(n370), .Z(n271) );
  GTECH_XOR2 U342 ( .A(n366), .B(n371), .Z(n370) );
  GTECH_NOT U343 ( .A(n372), .Z(n371) );
  GTECH_XOR2 U344 ( .A(n273), .B(n253), .Z(n366) );
  GTECH_OAI21 U345 ( .A(n12), .B(n369), .C(n373), .Z(N135) );
  GTECH_OAI21 U346 ( .A(n301), .B(n297), .C(n279), .Z(n373) );
  GTECH_OAI21 U347 ( .A(n12), .B(n374), .C(n368), .Z(n279) );
  GTECH_NOT U348 ( .A(n375), .Z(n297) );
  GTECH_NAND3 U349 ( .A(n28), .B(n376), .C(N155), .Z(n375) );
  GTECH_NOT U350 ( .A(n377), .Z(n301) );
  GTECH_NAND3 U351 ( .A(n10), .B(n378), .C(N155), .Z(n377) );
  GTECH_NAND2 U352 ( .A(n379), .B(N155), .Z(n369) );
  GTECH_XOR2 U353 ( .A(n376), .B(n28), .Z(n379) );
  GTECH_AND2 U354 ( .A(N155), .B(n380), .Z(N134) );
  GTECH_NOT U355 ( .A(n13), .Z(n380) );
  GTECH_AND2 U356 ( .A(N155), .B(n381), .Z(N133) );
  GTECH_NOT U357 ( .A(n14), .Z(n381) );
  GTECH_AND2 U358 ( .A(N155), .B(n382), .Z(N132) );
  GTECH_NOT U359 ( .A(n15), .Z(n382) );
  GTECH_AND2 U360 ( .A(N155), .B(n383), .Z(N131) );
  GTECH_NOT U361 ( .A(n16), .Z(n383) );
  GTECH_AND2 U362 ( .A(N155), .B(n384), .Z(N130) );
  GTECH_NOT U363 ( .A(n17), .Z(n384) );
  GTECH_AND2 U364 ( .A(N155), .B(n385), .Z(N129) );
  GTECH_NOT U365 ( .A(n18), .Z(n385) );
  GTECH_AND2 U366 ( .A(N155), .B(n386), .Z(N128) );
  GTECH_NOT U367 ( .A(n19), .Z(n386) );
  GTECH_AND2 U368 ( .A(N155), .B(n387), .Z(N127) );
  GTECH_NOT U369 ( .A(n20), .Z(n387) );
  GTECH_AND2 U370 ( .A(N155), .B(n388), .Z(N126) );
  GTECH_NOT U371 ( .A(n21), .Z(n388) );
  GTECH_AND2 U372 ( .A(N155), .B(n389), .Z(N125) );
  GTECH_NOT U373 ( .A(n22), .Z(n389) );
  GTECH_AND2 U374 ( .A(N155), .B(n390), .Z(N124) );
  GTECH_NOT U375 ( .A(n23), .Z(n390) );
  GTECH_AND2 U376 ( .A(N155), .B(n391), .Z(N123) );
  GTECH_NOT U377 ( .A(n24), .Z(n391) );
  GTECH_AND2 U378 ( .A(N155), .B(n392), .Z(N122) );
  GTECH_NOT U379 ( .A(n25), .Z(n392) );
  GTECH_AND2 U380 ( .A(N155), .B(n393), .Z(N121) );
  GTECH_NOT U381 ( .A(n26), .Z(n393) );
  GTECH_AND2 U382 ( .A(N155), .B(n394), .Z(N120) );
  GTECH_NOT U383 ( .A(n27), .Z(n394) );
  GTECH_NOT U384 ( .A(n303), .Z(N155) );
  GTECH_NAND4 U385 ( .A(n8), .B(n7), .C(n9), .D(n395), .Z(n303) );
  GTECH_AND3 U386 ( .A(n290), .B(n311), .C(n6), .Z(n395) );
  GTECH_NOT U387 ( .A(n251), .Z(n311) );
  GTECH_NOT U388 ( .A(n396), .Z(N116) );
  GTECH_AOI222 U389 ( .A(n272), .B(n300), .C(n274), .D(n302), .E(n298), .F(
        n270), .Z(n396) );
  GTECH_XOR2 U390 ( .A(n397), .B(n398), .Z(n298) );
  GTECH_ADD_ABC U391 ( .A(n31), .B(n267), .C(n399), .COUT(n398) );
  GTECH_XOR2 U392 ( .A(n400), .B(n397), .Z(n302) );
  GTECH_XOR2 U393 ( .A(A[16]), .B(n30), .Z(n397) );
  GTECH_OAI21 U394 ( .A(n401), .B(n31), .C(n402), .Z(n400) );
  GTECH_OAI21 U395 ( .A(n267), .B(n306), .C(n403), .Z(n402) );
  GTECH_NOT U396 ( .A(n30), .Z(n300) );
  GTECH_NAND2 U397 ( .A(n283), .B(n404), .Z(N115) );
  GTECH_NOT U398 ( .A(N41), .Z(n404) );
  GTECH_NAND2 U399 ( .A(n290), .B(n284), .Z(N41) );
  GTECH_NAND2 U400 ( .A(Ld), .B(n290), .Z(n284) );
  GTECH_NOT U401 ( .A(n405), .Z(N113) );
  GTECH_AOI222 U402 ( .A(n272), .B(n306), .C(n274), .D(n307), .E(n305), .F(
        n270), .Z(n405) );
  GTECH_XOR2 U403 ( .A(n406), .B(n399), .Z(n305) );
  GTECH_ADD_ABC U404 ( .A(n32), .B(n266), .C(n407), .COUT(n399) );
  GTECH_NOT U405 ( .A(n408), .Z(n307) );
  GTECH_XOR2 U406 ( .A(n406), .B(n409), .Z(n408) );
  GTECH_NOT U407 ( .A(n403), .Z(n409) );
  GTECH_OAI21 U408 ( .A(n32), .B(n410), .C(n411), .Z(n403) );
  GTECH_OAI21 U409 ( .A(n266), .B(n314), .C(n412), .Z(n411) );
  GTECH_XOR2 U410 ( .A(n401), .B(n31), .Z(n406) );
  GTECH_NOT U411 ( .A(n267), .Z(n401) );
  GTECH_NOT U412 ( .A(n31), .Z(n306) );
  GTECH_NOT U413 ( .A(n413), .Z(N112) );
  GTECH_AOI222 U414 ( .A(n272), .B(n314), .C(n274), .D(n315), .E(n313), .F(
        n270), .Z(n413) );
  GTECH_XOR2 U415 ( .A(n414), .B(n407), .Z(n313) );
  GTECH_ADD_ABC U416 ( .A(n33), .B(n265), .C(n415), .COUT(n407) );
  GTECH_NOT U417 ( .A(n416), .Z(n315) );
  GTECH_XOR2 U418 ( .A(n414), .B(n417), .Z(n416) );
  GTECH_NOT U419 ( .A(n412), .Z(n417) );
  GTECH_OAI21 U420 ( .A(n33), .B(n418), .C(n419), .Z(n412) );
  GTECH_OAI21 U421 ( .A(n265), .B(n318), .C(n420), .Z(n419) );
  GTECH_XOR2 U422 ( .A(n410), .B(n32), .Z(n414) );
  GTECH_NOT U423 ( .A(n266), .Z(n410) );
  GTECH_NOT U424 ( .A(n32), .Z(n314) );
  GTECH_NOT U425 ( .A(n421), .Z(N111) );
  GTECH_AOI222 U426 ( .A(n272), .B(n318), .C(n274), .D(n319), .E(n317), .F(
        n270), .Z(n421) );
  GTECH_XOR2 U427 ( .A(n422), .B(n415), .Z(n317) );
  GTECH_ADD_ABC U428 ( .A(n34), .B(n264), .C(n423), .COUT(n415) );
  GTECH_NOT U429 ( .A(n424), .Z(n319) );
  GTECH_XOR2 U430 ( .A(n422), .B(n425), .Z(n424) );
  GTECH_NOT U431 ( .A(n420), .Z(n425) );
  GTECH_OAI21 U432 ( .A(n34), .B(n426), .C(n427), .Z(n420) );
  GTECH_OAI21 U433 ( .A(n264), .B(n322), .C(n428), .Z(n427) );
  GTECH_XOR2 U434 ( .A(n418), .B(n33), .Z(n422) );
  GTECH_NOT U435 ( .A(n265), .Z(n418) );
  GTECH_NOT U436 ( .A(n33), .Z(n318) );
  GTECH_NOT U437 ( .A(n429), .Z(N110) );
  GTECH_AOI222 U438 ( .A(n272), .B(n322), .C(n274), .D(n323), .E(n321), .F(
        n270), .Z(n429) );
  GTECH_XOR2 U439 ( .A(n430), .B(n423), .Z(n321) );
  GTECH_ADD_ABC U440 ( .A(n35), .B(n263), .C(n431), .COUT(n423) );
  GTECH_NOT U441 ( .A(n432), .Z(n323) );
  GTECH_XOR2 U442 ( .A(n430), .B(n433), .Z(n432) );
  GTECH_NOT U443 ( .A(n428), .Z(n433) );
  GTECH_OAI21 U444 ( .A(n35), .B(n434), .C(n435), .Z(n428) );
  GTECH_OAI21 U445 ( .A(n263), .B(n326), .C(n436), .Z(n435) );
  GTECH_XOR2 U446 ( .A(n426), .B(n34), .Z(n430) );
  GTECH_NOT U447 ( .A(n264), .Z(n426) );
  GTECH_NOT U448 ( .A(n34), .Z(n322) );
  GTECH_NOT U449 ( .A(n437), .Z(N109) );
  GTECH_AOI222 U450 ( .A(n272), .B(n326), .C(n274), .D(n327), .E(n325), .F(
        n270), .Z(n437) );
  GTECH_XOR2 U451 ( .A(n438), .B(n431), .Z(n325) );
  GTECH_ADD_ABC U452 ( .A(n36), .B(n262), .C(n439), .COUT(n431) );
  GTECH_NOT U453 ( .A(n440), .Z(n327) );
  GTECH_XOR2 U454 ( .A(n438), .B(n441), .Z(n440) );
  GTECH_NOT U455 ( .A(n436), .Z(n441) );
  GTECH_OAI21 U456 ( .A(n36), .B(n442), .C(n443), .Z(n436) );
  GTECH_OAI21 U457 ( .A(n262), .B(n330), .C(n444), .Z(n443) );
  GTECH_XOR2 U458 ( .A(n434), .B(n35), .Z(n438) );
  GTECH_NOT U459 ( .A(n263), .Z(n434) );
  GTECH_NOT U460 ( .A(n35), .Z(n326) );
  GTECH_NOT U461 ( .A(n445), .Z(N108) );
  GTECH_AOI222 U462 ( .A(n272), .B(n330), .C(n274), .D(n331), .E(n329), .F(
        n270), .Z(n445) );
  GTECH_XOR2 U463 ( .A(n446), .B(n439), .Z(n329) );
  GTECH_ADD_ABC U464 ( .A(n37), .B(n261), .C(n447), .COUT(n439) );
  GTECH_NOT U465 ( .A(n448), .Z(n331) );
  GTECH_XOR2 U466 ( .A(n446), .B(n449), .Z(n448) );
  GTECH_NOT U467 ( .A(n444), .Z(n449) );
  GTECH_OAI21 U468 ( .A(n37), .B(n450), .C(n451), .Z(n444) );
  GTECH_OAI21 U469 ( .A(n261), .B(n334), .C(n452), .Z(n451) );
  GTECH_XOR2 U470 ( .A(n442), .B(n36), .Z(n446) );
  GTECH_NOT U471 ( .A(n262), .Z(n442) );
  GTECH_NOT U472 ( .A(n36), .Z(n330) );
  GTECH_NOT U473 ( .A(n453), .Z(N107) );
  GTECH_AOI222 U474 ( .A(n272), .B(n334), .C(n274), .D(n335), .E(n333), .F(
        n270), .Z(n453) );
  GTECH_XOR2 U475 ( .A(n454), .B(n447), .Z(n333) );
  GTECH_ADD_ABC U476 ( .A(n38), .B(n260), .C(n455), .COUT(n447) );
  GTECH_NOT U477 ( .A(n456), .Z(n335) );
  GTECH_XOR2 U478 ( .A(n454), .B(n457), .Z(n456) );
  GTECH_NOT U479 ( .A(n452), .Z(n457) );
  GTECH_OAI21 U480 ( .A(n38), .B(n458), .C(n459), .Z(n452) );
  GTECH_OAI21 U481 ( .A(n260), .B(n338), .C(n460), .Z(n459) );
  GTECH_XOR2 U482 ( .A(n450), .B(n37), .Z(n454) );
  GTECH_NOT U483 ( .A(n261), .Z(n450) );
  GTECH_NOT U484 ( .A(n37), .Z(n334) );
  GTECH_NOT U485 ( .A(n461), .Z(N106) );
  GTECH_AOI222 U486 ( .A(n272), .B(n338), .C(n274), .D(n339), .E(n337), .F(
        n270), .Z(n461) );
  GTECH_XOR2 U487 ( .A(n462), .B(n455), .Z(n337) );
  GTECH_ADD_ABC U488 ( .A(n39), .B(n259), .C(n463), .COUT(n455) );
  GTECH_NOT U489 ( .A(n464), .Z(n339) );
  GTECH_XOR2 U490 ( .A(n462), .B(n465), .Z(n464) );
  GTECH_NOT U491 ( .A(n460), .Z(n465) );
  GTECH_OAI21 U492 ( .A(n39), .B(n466), .C(n467), .Z(n460) );
  GTECH_OAI21 U493 ( .A(n259), .B(n342), .C(n468), .Z(n467) );
  GTECH_XOR2 U494 ( .A(n458), .B(n38), .Z(n462) );
  GTECH_NOT U495 ( .A(n260), .Z(n458) );
  GTECH_NOT U496 ( .A(n38), .Z(n338) );
  GTECH_NOT U497 ( .A(n469), .Z(N105) );
  GTECH_AOI222 U498 ( .A(n272), .B(n342), .C(n274), .D(n343), .E(n341), .F(
        n270), .Z(n469) );
  GTECH_XOR2 U499 ( .A(n470), .B(n463), .Z(n341) );
  GTECH_ADD_ABC U500 ( .A(n40), .B(n258), .C(n471), .COUT(n463) );
  GTECH_NOT U501 ( .A(n472), .Z(n343) );
  GTECH_XOR2 U502 ( .A(n470), .B(n473), .Z(n472) );
  GTECH_NOT U503 ( .A(n468), .Z(n473) );
  GTECH_OAI21 U504 ( .A(n40), .B(n474), .C(n475), .Z(n468) );
  GTECH_OAI21 U505 ( .A(n258), .B(n346), .C(n476), .Z(n475) );
  GTECH_XOR2 U506 ( .A(n466), .B(n39), .Z(n470) );
  GTECH_NOT U507 ( .A(n259), .Z(n466) );
  GTECH_NOT U508 ( .A(n39), .Z(n342) );
  GTECH_NOT U509 ( .A(n477), .Z(N104) );
  GTECH_AOI222 U510 ( .A(n272), .B(n346), .C(n274), .D(n347), .E(n345), .F(
        n270), .Z(n477) );
  GTECH_XOR2 U511 ( .A(n478), .B(n471), .Z(n345) );
  GTECH_ADD_ABC U512 ( .A(n41), .B(n257), .C(n479), .COUT(n471) );
  GTECH_NOT U513 ( .A(n480), .Z(n347) );
  GTECH_XOR2 U514 ( .A(n478), .B(n481), .Z(n480) );
  GTECH_NOT U515 ( .A(n476), .Z(n481) );
  GTECH_OAI21 U516 ( .A(n41), .B(n482), .C(n483), .Z(n476) );
  GTECH_OAI21 U517 ( .A(n257), .B(n350), .C(n484), .Z(n483) );
  GTECH_XOR2 U518 ( .A(n474), .B(n40), .Z(n478) );
  GTECH_NOT U519 ( .A(n258), .Z(n474) );
  GTECH_NOT U520 ( .A(n40), .Z(n346) );
  GTECH_NOT U521 ( .A(n485), .Z(N103) );
  GTECH_AOI222 U522 ( .A(n272), .B(n350), .C(n274), .D(n351), .E(n349), .F(
        n270), .Z(n485) );
  GTECH_XOR2 U523 ( .A(n486), .B(n479), .Z(n349) );
  GTECH_ADD_ABC U524 ( .A(n42), .B(n256), .C(n487), .COUT(n479) );
  GTECH_NOT U525 ( .A(n488), .Z(n351) );
  GTECH_XOR2 U526 ( .A(n486), .B(n489), .Z(n488) );
  GTECH_NOT U527 ( .A(n484), .Z(n489) );
  GTECH_OAI21 U528 ( .A(n42), .B(n490), .C(n491), .Z(n484) );
  GTECH_OAI21 U529 ( .A(n256), .B(n354), .C(n492), .Z(n491) );
  GTECH_XOR2 U530 ( .A(n482), .B(n41), .Z(n486) );
  GTECH_NOT U531 ( .A(n257), .Z(n482) );
  GTECH_NOT U532 ( .A(n41), .Z(n350) );
  GTECH_NOT U533 ( .A(n493), .Z(N102) );
  GTECH_AOI222 U534 ( .A(n272), .B(n354), .C(n274), .D(n355), .E(n353), .F(
        n270), .Z(n493) );
  GTECH_XOR2 U535 ( .A(n494), .B(n487), .Z(n353) );
  GTECH_ADD_ABC U536 ( .A(n43), .B(n255), .C(n495), .COUT(n487) );
  GTECH_NOT U537 ( .A(n496), .Z(n355) );
  GTECH_XOR2 U538 ( .A(n494), .B(n497), .Z(n496) );
  GTECH_NOT U539 ( .A(n492), .Z(n497) );
  GTECH_OAI21 U540 ( .A(n43), .B(n498), .C(n499), .Z(n492) );
  GTECH_OAI21 U541 ( .A(n255), .B(n358), .C(n500), .Z(n499) );
  GTECH_XOR2 U542 ( .A(n490), .B(n42), .Z(n494) );
  GTECH_NOT U543 ( .A(n256), .Z(n490) );
  GTECH_NOT U544 ( .A(n42), .Z(n354) );
  GTECH_NOT U545 ( .A(n501), .Z(N101) );
  GTECH_AOI222 U546 ( .A(n272), .B(n358), .C(n274), .D(n359), .E(n357), .F(
        n270), .Z(n501) );
  GTECH_XOR2 U547 ( .A(n502), .B(n495), .Z(n357) );
  GTECH_ADD_ABC U548 ( .A(n29), .B(n254), .C(n503), .COUT(n495) );
  GTECH_NOT U549 ( .A(n504), .Z(n359) );
  GTECH_XOR2 U550 ( .A(n502), .B(n505), .Z(n504) );
  GTECH_NOT U551 ( .A(n500), .Z(n505) );
  GTECH_OAI21 U552 ( .A(n29), .B(n506), .C(n507), .Z(n500) );
  GTECH_OAI21 U553 ( .A(n254), .B(n362), .C(n508), .Z(n507) );
  GTECH_XOR2 U554 ( .A(n498), .B(n43), .Z(n502) );
  GTECH_NOT U555 ( .A(n255), .Z(n498) );
  GTECH_NOT U556 ( .A(n43), .Z(n358) );
  GTECH_NOT U557 ( .A(n509), .Z(N100) );
  GTECH_AOI222 U558 ( .A(n361), .B(n270), .C(n272), .D(n362), .E(n274), .F(
        n363), .Z(n509) );
  GTECH_NOT U559 ( .A(n510), .Z(n363) );
  GTECH_XOR2 U560 ( .A(n511), .B(n512), .Z(n510) );
  GTECH_NOT U561 ( .A(n508), .Z(n512) );
  GTECH_OAI21 U562 ( .A(n11), .B(n513), .C(n514), .Z(n508) );
  GTECH_OAI21 U563 ( .A(n253), .B(n273), .C(n368), .Z(n514) );
  GTECH_NAND2 U564 ( .A(n12), .B(n374), .Z(n368) );
  GTECH_NOT U565 ( .A(n11), .Z(n273) );
  GTECH_NOT U566 ( .A(n253), .Z(n513) );
  GTECH_NOT U567 ( .A(n282), .Z(n274) );
  GTECH_NAND2 U568 ( .A(N82), .B(n10), .Z(n282) );
  GTECH_NOT U569 ( .A(n515), .Z(N82) );
  GTECH_NOT U570 ( .A(n29), .Z(n362) );
  GTECH_OAI21 U571 ( .A(n10), .B(n515), .C(n516), .Z(n272) );
  GTECH_NAND3 U572 ( .A(n28), .B(n288), .C(n10), .Z(n516) );
  GTECH_NAND2 U573 ( .A(n288), .B(n378), .Z(n515) );
  GTECH_NOT U574 ( .A(n28), .Z(n378) );
  GTECH_NOT U575 ( .A(n281), .Z(n270) );
  GTECH_NAND3 U576 ( .A(n288), .B(n376), .C(n28), .Z(n281) );
  GTECH_NOT U577 ( .A(n10), .Z(n376) );
  GTECH_NOT U578 ( .A(n283), .Z(n288) );
  GTECH_OAI21 U579 ( .A(n286), .B(n287), .C(n517), .Z(n283) );
  GTECH_AND2 U580 ( .A(n289), .B(n290), .Z(n517) );
  GTECH_NOT U581 ( .A(Rst), .Z(n290) );
  GTECH_NOT U582 ( .A(Ld), .Z(n289) );
  GTECH_NOT U583 ( .A(n9), .Z(n287) );
  GTECH_NAND2 U584 ( .A(n8), .B(n292), .Z(n286) );
  GTECH_NOT U585 ( .A(n295), .Z(n292) );
  GTECH_NAND2 U586 ( .A(n7), .B(n294), .Z(n295) );
  GTECH_NOT U587 ( .A(n518), .Z(n294) );
  GTECH_NAND2 U588 ( .A(n6), .B(n251), .Z(n518) );
  GTECH_XOR2 U589 ( .A(n511), .B(n503), .Z(n361) );
  GTECH_ADD_ABC U590 ( .A(n253), .B(n11), .C(n372), .COUT(n503) );
  GTECH_NAND2 U591 ( .A(n277), .B(n374), .Z(n372) );
  GTECH_NOT U592 ( .A(n252), .Z(n374) );
  GTECH_NOT U593 ( .A(n12), .Z(n277) );
  GTECH_XOR2 U594 ( .A(n506), .B(n29), .Z(n511) );
  GTECH_NOT U595 ( .A(n254), .Z(n506) );
endmodule

