
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_XOR2 U75 ( .A(n83), .B(n84), .Z(N155) );
  GTECH_AND2 U76 ( .A(n85), .B(n86), .Z(n84) );
  GTECH_OAI22 U77 ( .A(n87), .B(n88), .C(n89), .D(n90), .Z(n83) );
  GTECH_NOT U78 ( .A(n91), .Z(n90) );
  GTECH_XOR2 U79 ( .A(n85), .B(n86), .Z(N154) );
  GTECH_NOT U80 ( .A(n92), .Z(n86) );
  GTECH_XOR2 U81 ( .A(n91), .B(n89), .Z(n92) );
  GTECH_AOI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n89) );
  GTECH_NAND2 U83 ( .A(n95), .B(n96), .Z(n94) );
  GTECH_XOR2 U84 ( .A(n88), .B(n87), .Z(n91) );
  GTECH_OA22 U85 ( .A(n97), .B(n98), .C(n99), .D(n100), .Z(n87) );
  GTECH_AND2 U86 ( .A(n97), .B(n98), .Z(n99) );
  GTECH_NAND2 U87 ( .A(I_b[7]), .B(I_a[7]), .Z(n88) );
  GTECH_NOT U88 ( .A(n101), .Z(n85) );
  GTECH_NAND2 U89 ( .A(n102), .B(n103), .Z(n101) );
  GTECH_XOR2 U90 ( .A(n102), .B(n103), .Z(N153) );
  GTECH_NOT U91 ( .A(n104), .Z(n103) );
  GTECH_NAND2 U92 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_XOR3 U93 ( .A(n107), .B(n108), .C(n95), .Z(n102) );
  GTECH_XOR3 U94 ( .A(n109), .B(n110), .C(n100), .Z(n95) );
  GTECH_OAI22 U95 ( .A(n111), .B(n112), .C(n113), .D(n114), .Z(n100) );
  GTECH_NOR2 U96 ( .A(n115), .B(n116), .Z(n111) );
  GTECH_NOT U97 ( .A(n98), .Z(n110) );
  GTECH_NAND2 U98 ( .A(I_a[7]), .B(I_b[6]), .Z(n98) );
  GTECH_NOT U99 ( .A(n97), .Z(n109) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n97) );
  GTECH_NOT U101 ( .A(n93), .Z(n108) );
  GTECH_AO22 U102 ( .A(n117), .B(n118), .C(n119), .D(n120), .Z(n93) );
  GTECH_OR2 U103 ( .A(n120), .B(n119), .Z(n118) );
  GTECH_NOT U104 ( .A(n96), .Z(n107) );
  GTECH_NAND2 U105 ( .A(I_a[7]), .B(n121), .Z(n96) );
  GTECH_XOR2 U106 ( .A(n122), .B(n123), .Z(N152) );
  GTECH_NOT U107 ( .A(n105), .Z(n123) );
  GTECH_XOR3 U108 ( .A(n124), .B(n125), .C(n119), .Z(n105) );
  GTECH_XOR2 U109 ( .A(n126), .B(n121), .Z(n119) );
  GTECH_OAI21 U110 ( .A(n127), .B(n128), .C(n129), .Z(n121) );
  GTECH_AO21 U111 ( .A(n127), .B(n128), .C(n130), .Z(n129) );
  GTECH_AND2 U112 ( .A(I_a[7]), .B(I_b[5]), .Z(n126) );
  GTECH_NOT U113 ( .A(n120), .Z(n125) );
  GTECH_XOR3 U114 ( .A(n113), .B(n114), .C(n112), .Z(n120) );
  GTECH_OAI21 U115 ( .A(n131), .B(n132), .C(n133), .Z(n112) );
  GTECH_OAI21 U116 ( .A(n134), .B(n135), .C(n136), .Z(n133) );
  GTECH_NOT U117 ( .A(n116), .Z(n114) );
  GTECH_NAND2 U118 ( .A(I_b[6]), .B(I_a[6]), .Z(n116) );
  GTECH_NOT U119 ( .A(n115), .Z(n113) );
  GTECH_NAND2 U120 ( .A(I_b[7]), .B(I_a[5]), .Z(n115) );
  GTECH_NOT U121 ( .A(n117), .Z(n124) );
  GTECH_OAI2N2 U122 ( .A(n137), .B(n138), .C(n139), .D(n140), .Z(n117) );
  GTECH_OR_NOT U123 ( .A(n141), .B(n137), .Z(n140) );
  GTECH_NOT U124 ( .A(n106), .Z(n122) );
  GTECH_OAI21 U125 ( .A(n142), .B(n143), .C(n144), .Z(n106) );
  GTECH_OAI21 U126 ( .A(n145), .B(n146), .C(n147), .Z(n144) );
  GTECH_XOR3 U127 ( .A(n148), .B(n142), .C(n145), .Z(N151) );
  GTECH_NOT U128 ( .A(n143), .Z(n145) );
  GTECH_XOR3 U129 ( .A(n149), .B(n138), .C(n137), .Z(n143) );
  GTECH_XOR3 U130 ( .A(n150), .B(n151), .C(n130), .Z(n137) );
  GTECH_OAI22 U131 ( .A(n152), .B(n153), .C(n154), .D(n155), .Z(n130) );
  GTECH_NOR2 U132 ( .A(n156), .B(n157), .Z(n152) );
  GTECH_NOT U133 ( .A(n128), .Z(n151) );
  GTECH_NAND2 U134 ( .A(I_a[7]), .B(I_b[4]), .Z(n128) );
  GTECH_NOT U135 ( .A(n127), .Z(n150) );
  GTECH_NAND2 U136 ( .A(I_a[6]), .B(I_b[5]), .Z(n127) );
  GTECH_NOT U137 ( .A(n141), .Z(n138) );
  GTECH_XOR3 U138 ( .A(n135), .B(n134), .C(n136), .Z(n141) );
  GTECH_OAI21 U139 ( .A(n158), .B(n159), .C(n160), .Z(n136) );
  GTECH_OAI21 U140 ( .A(n161), .B(n162), .C(n163), .Z(n160) );
  GTECH_NOT U141 ( .A(n132), .Z(n134) );
  GTECH_NAND2 U142 ( .A(I_b[6]), .B(I_a[5]), .Z(n132) );
  GTECH_NOT U143 ( .A(n131), .Z(n135) );
  GTECH_NAND2 U144 ( .A(I_b[7]), .B(I_a[4]), .Z(n131) );
  GTECH_NOT U145 ( .A(n139), .Z(n149) );
  GTECH_AO22 U146 ( .A(n164), .B(n165), .C(n166), .D(n167), .Z(n139) );
  GTECH_OR2 U147 ( .A(n167), .B(n166), .Z(n165) );
  GTECH_NOT U148 ( .A(n146), .Z(n142) );
  GTECH_OAI22 U149 ( .A(n168), .B(n169), .C(n170), .D(n171), .Z(n146) );
  GTECH_NOT U150 ( .A(I_a[7]), .Z(n171) );
  GTECH_NOT U151 ( .A(n172), .Z(n169) );
  GTECH_NOT U152 ( .A(n147), .Z(n148) );
  GTECH_OAI21 U153 ( .A(n173), .B(n174), .C(n175), .Z(n147) );
  GTECH_OAI21 U154 ( .A(n176), .B(n177), .C(n178), .Z(n175) );
  GTECH_XOR3 U155 ( .A(n179), .B(n174), .C(n177), .Z(N150) );
  GTECH_NOT U156 ( .A(n173), .Z(n177) );
  GTECH_XOR2 U157 ( .A(n172), .B(n168), .Z(n173) );
  GTECH_AND2 U158 ( .A(n180), .B(n181), .Z(n168) );
  GTECH_OR_NOT U159 ( .A(n182), .B(n183), .Z(n181) );
  GTECH_OAI21 U160 ( .A(n184), .B(n183), .C(n185), .Z(n180) );
  GTECH_XOR2 U161 ( .A(n186), .B(n170), .Z(n172) );
  GTECH_AOI2N2 U162 ( .A(n187), .B(n188), .C(n189), .D(n190), .Z(n170) );
  GTECH_NAND2 U163 ( .A(n189), .B(n190), .Z(n188) );
  GTECH_NAND2 U164 ( .A(I_a[7]), .B(I_b[3]), .Z(n186) );
  GTECH_NOT U165 ( .A(n176), .Z(n174) );
  GTECH_XOR3 U166 ( .A(n191), .B(n192), .C(n166), .Z(n176) );
  GTECH_XOR3 U167 ( .A(n154), .B(n155), .C(n153), .Z(n166) );
  GTECH_OAI21 U168 ( .A(n193), .B(n194), .C(n195), .Z(n153) );
  GTECH_OAI21 U169 ( .A(n196), .B(n197), .C(n198), .Z(n195) );
  GTECH_NOT U170 ( .A(n157), .Z(n155) );
  GTECH_NAND2 U171 ( .A(I_a[6]), .B(I_b[4]), .Z(n157) );
  GTECH_NOT U172 ( .A(n156), .Z(n154) );
  GTECH_NAND2 U173 ( .A(I_b[5]), .B(I_a[5]), .Z(n156) );
  GTECH_NOT U174 ( .A(n167), .Z(n192) );
  GTECH_XOR3 U175 ( .A(n162), .B(n161), .C(n163), .Z(n167) );
  GTECH_OAI21 U176 ( .A(n199), .B(n200), .C(n201), .Z(n163) );
  GTECH_OAI21 U177 ( .A(n202), .B(n203), .C(n204), .Z(n201) );
  GTECH_NOT U178 ( .A(n159), .Z(n161) );
  GTECH_NAND2 U179 ( .A(I_b[6]), .B(I_a[4]), .Z(n159) );
  GTECH_NOT U180 ( .A(n158), .Z(n162) );
  GTECH_NAND2 U181 ( .A(I_b[7]), .B(I_a[3]), .Z(n158) );
  GTECH_NOT U182 ( .A(n164), .Z(n191) );
  GTECH_AO22 U183 ( .A(n205), .B(n206), .C(n207), .D(n208), .Z(n164) );
  GTECH_OR2 U184 ( .A(n208), .B(n207), .Z(n206) );
  GTECH_NOT U185 ( .A(n178), .Z(n179) );
  GTECH_OAI21 U186 ( .A(n209), .B(n210), .C(n211), .Z(n178) );
  GTECH_OAI21 U187 ( .A(n212), .B(n213), .C(n214), .Z(n211) );
  GTECH_XOR3 U188 ( .A(n215), .B(n210), .C(n213), .Z(N149) );
  GTECH_NOT U189 ( .A(n209), .Z(n213) );
  GTECH_XOR3 U190 ( .A(n184), .B(n216), .C(n183), .Z(n209) );
  GTECH_XOR3 U191 ( .A(n217), .B(n218), .C(n187), .Z(n183) );
  GTECH_OAI21 U192 ( .A(n219), .B(n220), .C(n221), .Z(n187) );
  GTECH_AO21 U193 ( .A(n219), .B(n220), .C(n222), .Z(n221) );
  GTECH_NOT U194 ( .A(n190), .Z(n218) );
  GTECH_NAND2 U195 ( .A(I_a[7]), .B(I_b[2]), .Z(n190) );
  GTECH_NOT U196 ( .A(n189), .Z(n217) );
  GTECH_NAND2 U197 ( .A(I_a[6]), .B(I_b[3]), .Z(n189) );
  GTECH_NOT U198 ( .A(n185), .Z(n216) );
  GTECH_OAI21 U199 ( .A(n223), .B(n224), .C(n225), .Z(n185) );
  GTECH_OAI21 U200 ( .A(n226), .B(n227), .C(n228), .Z(n225) );
  GTECH_NOT U201 ( .A(n226), .Z(n224) );
  GTECH_NOT U202 ( .A(n182), .Z(n184) );
  GTECH_NAND2 U203 ( .A(I_a[7]), .B(n229), .Z(n182) );
  GTECH_NOT U204 ( .A(n212), .Z(n210) );
  GTECH_XOR3 U205 ( .A(n230), .B(n231), .C(n207), .Z(n212) );
  GTECH_XOR3 U206 ( .A(n197), .B(n196), .C(n198), .Z(n207) );
  GTECH_OAI21 U207 ( .A(n232), .B(n233), .C(n234), .Z(n198) );
  GTECH_OAI21 U208 ( .A(n235), .B(n236), .C(n237), .Z(n234) );
  GTECH_NOT U209 ( .A(n194), .Z(n196) );
  GTECH_NAND2 U210 ( .A(I_a[5]), .B(I_b[4]), .Z(n194) );
  GTECH_NOT U211 ( .A(n193), .Z(n197) );
  GTECH_NAND2 U212 ( .A(I_b[5]), .B(I_a[4]), .Z(n193) );
  GTECH_NOT U213 ( .A(n208), .Z(n231) );
  GTECH_XOR3 U214 ( .A(n203), .B(n202), .C(n204), .Z(n208) );
  GTECH_OAI21 U215 ( .A(n238), .B(n239), .C(n240), .Z(n204) );
  GTECH_NOT U216 ( .A(n200), .Z(n202) );
  GTECH_NAND2 U217 ( .A(I_b[6]), .B(I_a[3]), .Z(n200) );
  GTECH_NOT U218 ( .A(n199), .Z(n203) );
  GTECH_NAND2 U219 ( .A(I_b[7]), .B(I_a[2]), .Z(n199) );
  GTECH_NOT U220 ( .A(n205), .Z(n230) );
  GTECH_OAI2N2 U221 ( .A(n241), .B(n242), .C(n243), .D(n244), .Z(n205) );
  GTECH_OR_NOT U222 ( .A(n245), .B(n241), .Z(n244) );
  GTECH_NOT U223 ( .A(n214), .Z(n215) );
  GTECH_OAI2N2 U224 ( .A(n246), .B(n247), .C(n248), .D(n249), .Z(n214) );
  GTECH_NAND2 U225 ( .A(n246), .B(n247), .Z(n249) );
  GTECH_XOR3 U226 ( .A(n250), .B(n251), .C(n246), .Z(N148) );
  GTECH_XOR3 U227 ( .A(n252), .B(n227), .C(n226), .Z(n246) );
  GTECH_XOR2 U228 ( .A(n253), .B(n229), .Z(n226) );
  GTECH_OAI21 U229 ( .A(n254), .B(n255), .C(n256), .Z(n229) );
  GTECH_AO21 U230 ( .A(n254), .B(n255), .C(n257), .Z(n256) );
  GTECH_AND2 U231 ( .A(I_a[7]), .B(I_b[1]), .Z(n253) );
  GTECH_NOT U232 ( .A(n223), .Z(n227) );
  GTECH_XOR3 U233 ( .A(n258), .B(n259), .C(n222), .Z(n223) );
  GTECH_OAI22 U234 ( .A(n260), .B(n261), .C(n262), .D(n263), .Z(n222) );
  GTECH_NOR2 U235 ( .A(n264), .B(n265), .Z(n260) );
  GTECH_NOT U236 ( .A(n220), .Z(n259) );
  GTECH_NAND2 U237 ( .A(I_a[6]), .B(I_b[2]), .Z(n220) );
  GTECH_NOT U238 ( .A(n219), .Z(n258) );
  GTECH_NAND2 U239 ( .A(I_a[5]), .B(I_b[3]), .Z(n219) );
  GTECH_NOT U240 ( .A(n228), .Z(n252) );
  GTECH_OAI21 U241 ( .A(n266), .B(n267), .C(n268), .Z(n228) );
  GTECH_OAI21 U242 ( .A(n269), .B(n270), .C(n271), .Z(n268) );
  GTECH_NOT U243 ( .A(n269), .Z(n267) );
  GTECH_NOT U244 ( .A(n247), .Z(n251) );
  GTECH_XOR3 U245 ( .A(n272), .B(n242), .C(n241), .Z(n247) );
  GTECH_XOR3 U246 ( .A(n273), .B(n274), .C(n240), .Z(n241) );
  GTECH_NAND3 U247 ( .A(I_b[6]), .B(I_a[1]), .C(n275), .Z(n240) );
  GTECH_NOT U248 ( .A(n239), .Z(n274) );
  GTECH_NAND2 U249 ( .A(I_b[6]), .B(I_a[2]), .Z(n239) );
  GTECH_NOT U250 ( .A(n238), .Z(n273) );
  GTECH_NAND2 U251 ( .A(I_b[7]), .B(I_a[1]), .Z(n238) );
  GTECH_NOT U252 ( .A(n245), .Z(n242) );
  GTECH_XOR3 U253 ( .A(n236), .B(n235), .C(n237), .Z(n245) );
  GTECH_OAI21 U254 ( .A(n276), .B(n277), .C(n278), .Z(n237) );
  GTECH_OAI21 U255 ( .A(n279), .B(n280), .C(n281), .Z(n278) );
  GTECH_NOT U256 ( .A(n233), .Z(n235) );
  GTECH_NAND2 U257 ( .A(I_a[4]), .B(I_b[4]), .Z(n233) );
  GTECH_NOT U258 ( .A(n232), .Z(n236) );
  GTECH_NAND2 U259 ( .A(I_b[5]), .B(I_a[3]), .Z(n232) );
  GTECH_NOT U260 ( .A(n243), .Z(n272) );
  GTECH_OAI22 U261 ( .A(n282), .B(n283), .C(n284), .D(n285), .Z(n243) );
  GTECH_AND_NOT U262 ( .A(n284), .B(n286), .Z(n282) );
  GTECH_NOT U263 ( .A(n248), .Z(n250) );
  GTECH_AO22 U264 ( .A(n287), .B(n288), .C(n289), .D(n290), .Z(n248) );
  GTECH_OR2 U265 ( .A(n290), .B(n289), .Z(n288) );
  GTECH_XOR3 U266 ( .A(n291), .B(n292), .C(n289), .Z(N147) );
  GTECH_XOR3 U267 ( .A(n293), .B(n285), .C(n284), .Z(n289) );
  GTECH_XOR2 U268 ( .A(n294), .B(n275), .Z(n284) );
  GTECH_NOT U269 ( .A(n295), .Z(n275) );
  GTECH_NAND2 U270 ( .A(I_b[7]), .B(I_a[0]), .Z(n295) );
  GTECH_NAND2 U271 ( .A(I_b[6]), .B(I_a[1]), .Z(n294) );
  GTECH_NOT U272 ( .A(n286), .Z(n285) );
  GTECH_XOR3 U273 ( .A(n280), .B(n279), .C(n281), .Z(n286) );
  GTECH_OAI21 U274 ( .A(n296), .B(n297), .C(n298), .Z(n281) );
  GTECH_NOT U275 ( .A(n277), .Z(n279) );
  GTECH_NAND2 U276 ( .A(I_a[3]), .B(I_b[4]), .Z(n277) );
  GTECH_NOT U277 ( .A(n276), .Z(n280) );
  GTECH_NAND2 U278 ( .A(I_b[5]), .B(I_a[2]), .Z(n276) );
  GTECH_NOT U279 ( .A(n283), .Z(n293) );
  GTECH_NAND2 U280 ( .A(n299), .B(n300), .Z(n283) );
  GTECH_NOT U281 ( .A(n301), .Z(n300) );
  GTECH_NOT U282 ( .A(n290), .Z(n292) );
  GTECH_XOR3 U283 ( .A(n271), .B(n270), .C(n269), .Z(n290) );
  GTECH_XOR3 U284 ( .A(n262), .B(n263), .C(n261), .Z(n269) );
  GTECH_OAI21 U285 ( .A(n302), .B(n303), .C(n304), .Z(n261) );
  GTECH_AO21 U286 ( .A(n302), .B(n303), .C(n305), .Z(n304) );
  GTECH_NOT U287 ( .A(n265), .Z(n263) );
  GTECH_NAND2 U288 ( .A(I_a[5]), .B(I_b[2]), .Z(n265) );
  GTECH_NOT U289 ( .A(n264), .Z(n262) );
  GTECH_NAND2 U290 ( .A(I_a[4]), .B(I_b[3]), .Z(n264) );
  GTECH_NOT U291 ( .A(n266), .Z(n270) );
  GTECH_XOR3 U292 ( .A(n306), .B(n307), .C(n257), .Z(n266) );
  GTECH_OAI22 U293 ( .A(n308), .B(n309), .C(n310), .D(n311), .Z(n257) );
  GTECH_NOR2 U294 ( .A(n312), .B(n313), .Z(n308) );
  GTECH_NOT U295 ( .A(n255), .Z(n307) );
  GTECH_NAND2 U296 ( .A(I_a[7]), .B(I_b[0]), .Z(n255) );
  GTECH_NOT U297 ( .A(n254), .Z(n306) );
  GTECH_NAND2 U298 ( .A(I_a[6]), .B(I_b[1]), .Z(n254) );
  GTECH_AOI2N2 U299 ( .A(n314), .B(n315), .C(n316), .D(n317), .Z(n271) );
  GTECH_OR_NOT U300 ( .A(n318), .B(n316), .Z(n315) );
  GTECH_NOT U301 ( .A(n287), .Z(n291) );
  GTECH_OAI2N2 U302 ( .A(n319), .B(n320), .C(n321), .D(n322), .Z(n287) );
  GTECH_NAND2 U303 ( .A(n319), .B(n320), .Z(n322) );
  GTECH_XOR3 U304 ( .A(n323), .B(n324), .C(n319), .Z(N146) );
  GTECH_XOR3 U305 ( .A(n314), .B(n317), .C(n316), .Z(n319) );
  GTECH_XOR3 U306 ( .A(n310), .B(n311), .C(n309), .Z(n316) );
  GTECH_OAI21 U307 ( .A(n325), .B(n326), .C(n327), .Z(n309) );
  GTECH_OAI21 U308 ( .A(n328), .B(n329), .C(n330), .Z(n327) );
  GTECH_NOT U309 ( .A(n313), .Z(n311) );
  GTECH_NAND2 U310 ( .A(I_a[6]), .B(I_b[0]), .Z(n313) );
  GTECH_NOT U311 ( .A(n312), .Z(n310) );
  GTECH_NAND2 U312 ( .A(I_a[5]), .B(I_b[1]), .Z(n312) );
  GTECH_NOT U313 ( .A(n318), .Z(n317) );
  GTECH_XOR3 U314 ( .A(n331), .B(n332), .C(n305), .Z(n318) );
  GTECH_OAI22 U315 ( .A(n333), .B(n334), .C(n335), .D(n336), .Z(n305) );
  GTECH_NOR2 U316 ( .A(n337), .B(n338), .Z(n333) );
  GTECH_NOT U317 ( .A(n303), .Z(n332) );
  GTECH_NAND2 U318 ( .A(I_a[4]), .B(I_b[2]), .Z(n303) );
  GTECH_NOT U319 ( .A(n302), .Z(n331) );
  GTECH_NAND2 U320 ( .A(I_a[3]), .B(I_b[3]), .Z(n302) );
  GTECH_AOI22 U321 ( .A(n339), .B(n340), .C(n341), .D(n342), .Z(n314) );
  GTECH_OR2 U322 ( .A(n340), .B(n339), .Z(n342) );
  GTECH_NOT U323 ( .A(n320), .Z(n324) );
  GTECH_XOR2 U324 ( .A(n301), .B(n299), .Z(n320) );
  GTECH_NOT U325 ( .A(n343), .Z(n299) );
  GTECH_NAND2 U326 ( .A(I_b[6]), .B(I_a[0]), .Z(n343) );
  GTECH_XOR3 U327 ( .A(n344), .B(n345), .C(n298), .Z(n301) );
  GTECH_NAND3 U328 ( .A(I_a[1]), .B(I_b[4]), .C(n346), .Z(n298) );
  GTECH_NOT U329 ( .A(n297), .Z(n345) );
  GTECH_NAND2 U330 ( .A(I_a[2]), .B(I_b[4]), .Z(n297) );
  GTECH_NOT U331 ( .A(n296), .Z(n344) );
  GTECH_NAND2 U332 ( .A(I_b[5]), .B(I_a[1]), .Z(n296) );
  GTECH_NOT U333 ( .A(n321), .Z(n323) );
  GTECH_OAI21 U334 ( .A(n347), .B(n348), .C(n349), .Z(n321) );
  GTECH_OAI21 U335 ( .A(n350), .B(n351), .C(n352), .Z(n349) );
  GTECH_XOR3 U336 ( .A(n352), .B(n350), .C(n351), .Z(N145) );
  GTECH_NOT U337 ( .A(n347), .Z(n351) );
  GTECH_XOR3 U338 ( .A(n341), .B(n353), .C(n339), .Z(n347) );
  GTECH_XOR3 U339 ( .A(n335), .B(n336), .C(n334), .Z(n339) );
  GTECH_OAI21 U340 ( .A(n354), .B(n355), .C(n356), .Z(n334) );
  GTECH_NOT U341 ( .A(n338), .Z(n336) );
  GTECH_NAND2 U342 ( .A(I_a[3]), .B(I_b[2]), .Z(n338) );
  GTECH_NOT U343 ( .A(n337), .Z(n335) );
  GTECH_NAND2 U344 ( .A(I_a[2]), .B(I_b[3]), .Z(n337) );
  GTECH_NOT U345 ( .A(n340), .Z(n353) );
  GTECH_XOR3 U346 ( .A(n329), .B(n328), .C(n330), .Z(n340) );
  GTECH_OAI21 U347 ( .A(n357), .B(n358), .C(n359), .Z(n330) );
  GTECH_OAI21 U348 ( .A(n360), .B(n361), .C(n362), .Z(n359) );
  GTECH_NOT U349 ( .A(n326), .Z(n328) );
  GTECH_NAND2 U350 ( .A(I_a[5]), .B(I_b[0]), .Z(n326) );
  GTECH_NOT U351 ( .A(n325), .Z(n329) );
  GTECH_NAND2 U352 ( .A(I_a[4]), .B(I_b[1]), .Z(n325) );
  GTECH_AOI2N2 U353 ( .A(n363), .B(n364), .C(n365), .D(n366), .Z(n341) );
  GTECH_OR_NOT U354 ( .A(n367), .B(n365), .Z(n364) );
  GTECH_NOT U355 ( .A(n348), .Z(n350) );
  GTECH_XOR2 U356 ( .A(n368), .B(n346), .Z(n348) );
  GTECH_NOT U357 ( .A(n369), .Z(n346) );
  GTECH_NAND2 U358 ( .A(I_b[5]), .B(I_a[0]), .Z(n369) );
  GTECH_NAND2 U359 ( .A(I_a[1]), .B(I_b[4]), .Z(n368) );
  GTECH_NOT U360 ( .A(n370), .Z(n352) );
  GTECH_NAND2 U361 ( .A(n371), .B(n372), .Z(n370) );
  GTECH_XOR2 U362 ( .A(n371), .B(n372), .Z(N144) );
  GTECH_NOT U363 ( .A(n373), .Z(n372) );
  GTECH_XOR3 U364 ( .A(n363), .B(n366), .C(n365), .Z(n373) );
  GTECH_XOR3 U365 ( .A(n361), .B(n360), .C(n362), .Z(n365) );
  GTECH_OAI21 U366 ( .A(n374), .B(n375), .C(n376), .Z(n362) );
  GTECH_OAI21 U367 ( .A(n377), .B(n378), .C(n379), .Z(n376) );
  GTECH_NOT U368 ( .A(n358), .Z(n360) );
  GTECH_NAND2 U369 ( .A(I_a[4]), .B(I_b[0]), .Z(n358) );
  GTECH_NOT U370 ( .A(n357), .Z(n361) );
  GTECH_NAND2 U371 ( .A(I_a[3]), .B(I_b[1]), .Z(n357) );
  GTECH_NOT U372 ( .A(n367), .Z(n366) );
  GTECH_XOR3 U373 ( .A(n380), .B(n381), .C(n356), .Z(n367) );
  GTECH_NAND2 U374 ( .A(n382), .B(n383), .Z(n356) );
  GTECH_NOT U375 ( .A(n384), .Z(n383) );
  GTECH_NOT U376 ( .A(n355), .Z(n381) );
  GTECH_NAND2 U377 ( .A(I_a[2]), .B(I_b[2]), .Z(n355) );
  GTECH_NOT U378 ( .A(n354), .Z(n380) );
  GTECH_NAND2 U379 ( .A(I_a[1]), .B(I_b[3]), .Z(n354) );
  GTECH_OA22 U380 ( .A(n385), .B(n386), .C(n387), .D(n388), .Z(n363) );
  GTECH_AND_NOT U381 ( .A(n385), .B(n389), .Z(n387) );
  GTECH_NOT U382 ( .A(n390), .Z(n371) );
  GTECH_NAND2 U383 ( .A(I_b[4]), .B(I_a[0]), .Z(n390) );
  GTECH_XOR3 U384 ( .A(n391), .B(n386), .C(n385), .Z(N143) );
  GTECH_XOR2 U385 ( .A(n384), .B(n382), .Z(n385) );
  GTECH_NOT U386 ( .A(n392), .Z(n382) );
  GTECH_NAND2 U387 ( .A(I_b[3]), .B(I_a[0]), .Z(n392) );
  GTECH_NAND2 U388 ( .A(I_b[2]), .B(I_a[1]), .Z(n384) );
  GTECH_NOT U389 ( .A(n389), .Z(n386) );
  GTECH_XOR3 U390 ( .A(n378), .B(n377), .C(n379), .Z(n389) );
  GTECH_OAI21 U391 ( .A(n393), .B(n394), .C(n395), .Z(n379) );
  GTECH_NOT U392 ( .A(n375), .Z(n377) );
  GTECH_NAND2 U393 ( .A(I_a[3]), .B(I_b[0]), .Z(n375) );
  GTECH_NOT U394 ( .A(n374), .Z(n378) );
  GTECH_NAND2 U395 ( .A(I_b[1]), .B(I_a[2]), .Z(n374) );
  GTECH_NOT U396 ( .A(n388), .Z(n391) );
  GTECH_NAND2 U397 ( .A(n396), .B(n397), .Z(n388) );
  GTECH_XOR2 U398 ( .A(n396), .B(n397), .Z(N142) );
  GTECH_NOT U399 ( .A(n398), .Z(n397) );
  GTECH_XOR3 U400 ( .A(n399), .B(n400), .C(n395), .Z(n398) );
  GTECH_NAND3 U401 ( .A(n401), .B(I_a[1]), .C(I_b[0]), .Z(n395) );
  GTECH_NOT U402 ( .A(n394), .Z(n400) );
  GTECH_NAND2 U403 ( .A(I_b[0]), .B(I_a[2]), .Z(n394) );
  GTECH_NOT U404 ( .A(n393), .Z(n399) );
  GTECH_NAND2 U405 ( .A(I_b[1]), .B(I_a[1]), .Z(n393) );
  GTECH_NOT U406 ( .A(n402), .Z(n396) );
  GTECH_NAND2 U407 ( .A(I_b[2]), .B(I_a[0]), .Z(n402) );
  GTECH_XOR2 U408 ( .A(n401), .B(n403), .Z(N141) );
  GTECH_AND2 U409 ( .A(I_b[0]), .B(I_a[1]), .Z(n403) );
  GTECH_NOT U410 ( .A(n404), .Z(n401) );
  GTECH_NAND2 U411 ( .A(I_b[1]), .B(I_a[0]), .Z(n404) );
  GTECH_AND2 U412 ( .A(I_b[0]), .B(I_a[0]), .Z(N140) );
endmodule

