
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145;

  GTECH_XOR2 U89 ( .A(n70), .B(n71), .Z(sum[9]) );
  GTECH_XOR2 U90 ( .A(n72), .B(n73), .Z(sum[8]) );
  GTECH_XNOR2 U91 ( .A(n74), .B(n75), .Z(sum[7]) );
  GTECH_AOI21 U92 ( .A(n76), .B(n77), .C(n78), .Z(n75) );
  GTECH_XOR2 U93 ( .A(n77), .B(n76), .Z(sum[6]) );
  GTECH_AO22 U94 ( .A(b[5]), .B(a[5]), .C(n79), .D(n80), .Z(n76) );
  GTECH_XOR2 U95 ( .A(n80), .B(n79), .Z(sum[5]) );
  GTECH_OAI2N2 U96 ( .A(n81), .B(n82), .C(a[4]), .D(b[4]), .Z(n79) );
  GTECH_XNOR2 U97 ( .A(n83), .B(n81), .Z(sum[4]) );
  GTECH_XNOR2 U98 ( .A(n84), .B(n85), .Z(sum[3]) );
  GTECH_AOI21 U99 ( .A(n86), .B(n87), .C(n88), .Z(n85) );
  GTECH_XOR2 U100 ( .A(n87), .B(n86), .Z(sum[2]) );
  GTECH_AO22 U101 ( .A(b[1]), .B(a[1]), .C(n89), .D(n90), .Z(n86) );
  GTECH_XOR2 U102 ( .A(n90), .B(n89), .Z(sum[1]) );
  GTECH_AO22 U103 ( .A(n91), .B(cin), .C(a[0]), .D(b[0]), .Z(n89) );
  GTECH_XNOR2 U104 ( .A(n92), .B(n93), .Z(sum[15]) );
  GTECH_OAI21 U105 ( .A(n94), .B(n95), .C(n96), .Z(n92) );
  GTECH_XOR2 U106 ( .A(n94), .B(n95), .Z(sum[14]) );
  GTECH_AOI2N2 U107 ( .A(b[13]), .B(a[13]), .C(n97), .D(n98), .Z(n94) );
  GTECH_XOR2 U108 ( .A(n98), .B(n97), .Z(sum[13]) );
  GTECH_AOI21 U109 ( .A(cout), .B(n99), .C(n100), .Z(n97) );
  GTECH_XNOR2 U110 ( .A(n101), .B(cout), .Z(sum[12]) );
  GTECH_XNOR2 U111 ( .A(n102), .B(n103), .Z(sum[11]) );
  GTECH_AO21 U112 ( .A(n104), .B(n105), .C(n106), .Z(n102) );
  GTECH_XOR2 U113 ( .A(n105), .B(n104), .Z(sum[10]) );
  GTECH_AO21 U114 ( .A(n70), .B(n71), .C(n107), .Z(n104) );
  GTECH_AO21 U115 ( .A(n73), .B(n72), .C(n108), .Z(n70) );
  GTECH_XOR2 U116 ( .A(cin), .B(n91), .Z(sum[0]) );
  GTECH_OAI21 U117 ( .A(n109), .B(n110), .C(n111), .Z(cout) );
  GTECH_NOT U118 ( .A(n73), .Z(n109) );
  GTECH_OAI21 U119 ( .A(n81), .B(n112), .C(n113), .Z(n73) );
  GTECH_OA21 U120 ( .A(n114), .B(n115), .C(n116), .Z(n81) );
  GTECH_NOT U121 ( .A(cin), .Z(n115) );
  GTECH_NOR3 U122 ( .A(n112), .B(n114), .C(n110), .Z(Pm) );
  GTECH_NAND5 U123 ( .A(n87), .B(n90), .C(n84), .D(n117), .E(n91), .Z(n114) );
  GTECH_XOR2 U124 ( .A(a[0]), .B(b[0]), .Z(n91) );
  GTECH_OAI21 U125 ( .A(n118), .B(n110), .C(n111), .Z(Gm) );
  GTECH_OA21 U126 ( .A(n119), .B(n93), .C(n120), .Z(n111) );
  GTECH_OA21 U127 ( .A(n121), .B(n95), .C(n96), .Z(n119) );
  GTECH_AOI2N2 U128 ( .A(b[13]), .B(a[13]), .C(n98), .D(n122), .Z(n121) );
  GTECH_OR4 U129 ( .A(n101), .B(n93), .C(n95), .D(n98), .Z(n110) );
  GTECH_XNOR2 U130 ( .A(a[13]), .B(b[13]), .Z(n98) );
  GTECH_OAI21 U131 ( .A(b[14]), .B(a[14]), .C(n96), .Z(n95) );
  GTECH_OR_NOT U132 ( .A(n123), .B(b[14]), .Z(n96) );
  GTECH_NOT U133 ( .A(a[14]), .Z(n123) );
  GTECH_OAI21 U134 ( .A(b[15]), .B(a[15]), .C(n120), .Z(n93) );
  GTECH_NOT U135 ( .A(n124), .Z(n120) );
  GTECH_AND2 U136 ( .A(b[15]), .B(a[15]), .Z(n124) );
  GTECH_NOT U137 ( .A(n99), .Z(n101) );
  GTECH_OA21 U138 ( .A(b[12]), .B(a[12]), .C(n122), .Z(n99) );
  GTECH_NOT U139 ( .A(n100), .Z(n122) );
  GTECH_AND2 U140 ( .A(a[12]), .B(b[12]), .Z(n100) );
  GTECH_OA21 U141 ( .A(n116), .B(n112), .C(n113), .Z(n118) );
  GTECH_OA21 U142 ( .A(n125), .B(n103), .C(n126), .Z(n113) );
  GTECH_OA21 U143 ( .A(n127), .B(n128), .C(n129), .Z(n125) );
  GTECH_NOT U144 ( .A(n105), .Z(n128) );
  GTECH_AOI21 U145 ( .A(n71), .B(n108), .C(n107), .Z(n127) );
  GTECH_NAND4 U146 ( .A(n72), .B(n130), .C(n105), .D(n71), .Z(n112) );
  GTECH_OA21 U147 ( .A(b[9]), .B(a[9]), .C(n131), .Z(n71) );
  GTECH_NOT U148 ( .A(n107), .Z(n131) );
  GTECH_AND2 U149 ( .A(b[9]), .B(a[9]), .Z(n107) );
  GTECH_OA21 U150 ( .A(b[10]), .B(a[10]), .C(n129), .Z(n105) );
  GTECH_NOT U151 ( .A(n106), .Z(n129) );
  GTECH_AND2 U152 ( .A(a[10]), .B(b[10]), .Z(n106) );
  GTECH_NOT U153 ( .A(n103), .Z(n130) );
  GTECH_OAI21 U154 ( .A(b[11]), .B(a[11]), .C(n126), .Z(n103) );
  GTECH_NOT U155 ( .A(n132), .Z(n126) );
  GTECH_AND2 U156 ( .A(b[11]), .B(a[11]), .Z(n132) );
  GTECH_OA21 U157 ( .A(b[8]), .B(a[8]), .C(n133), .Z(n72) );
  GTECH_NOT U158 ( .A(n108), .Z(n133) );
  GTECH_AND2 U159 ( .A(b[8]), .B(a[8]), .Z(n108) );
  GTECH_AOI222 U160 ( .A(n117), .B(n134), .C(b[7]), .D(a[7]), .E(n74), .F(n135), .Z(n116) );
  GTECH_AO21 U161 ( .A(n136), .B(n77), .C(n78), .Z(n135) );
  GTECH_AND2 U162 ( .A(b[6]), .B(a[6]), .Z(n78) );
  GTECH_OAI21 U163 ( .A(n137), .B(n138), .C(n139), .Z(n136) );
  GTECH_NAND3 U164 ( .A(a[4]), .B(n80), .C(b[4]), .Z(n139) );
  GTECH_OAI2N2 U165 ( .A(n140), .B(n141), .C(b[3]), .D(a[3]), .Z(n134) );
  GTECH_NOT U166 ( .A(n84), .Z(n141) );
  GTECH_XOR2 U167 ( .A(a[3]), .B(b[3]), .Z(n84) );
  GTECH_AOI21 U168 ( .A(n142), .B(n87), .C(n88), .Z(n140) );
  GTECH_AND2 U169 ( .A(b[2]), .B(a[2]), .Z(n88) );
  GTECH_XOR2 U170 ( .A(a[2]), .B(b[2]), .Z(n87) );
  GTECH_OAI21 U171 ( .A(n143), .B(n144), .C(n145), .Z(n142) );
  GTECH_NAND3 U172 ( .A(a[0]), .B(n90), .C(b[0]), .Z(n145) );
  GTECH_XOR2 U173 ( .A(n144), .B(n143), .Z(n90) );
  GTECH_NOT U174 ( .A(a[1]), .Z(n144) );
  GTECH_NOT U175 ( .A(b[1]), .Z(n143) );
  GTECH_AND4 U176 ( .A(n83), .B(n80), .C(n77), .D(n74), .Z(n117) );
  GTECH_XOR2 U177 ( .A(a[7]), .B(b[7]), .Z(n74) );
  GTECH_XOR2 U178 ( .A(a[6]), .B(b[6]), .Z(n77) );
  GTECH_XOR2 U179 ( .A(n138), .B(n137), .Z(n80) );
  GTECH_NOT U180 ( .A(b[5]), .Z(n137) );
  GTECH_NOT U181 ( .A(a[5]), .Z(n138) );
  GTECH_NOT U182 ( .A(n82), .Z(n83) );
  GTECH_XNOR2 U183 ( .A(a[4]), .B(b[4]), .Z(n82) );
endmodule

