
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384;

  GTECH_MUX2 U132 ( .A(n271), .B(n272), .S(n273), .Z(sum[9]) );
  GTECH_XOR2 U133 ( .A(n274), .B(n275), .Z(n272) );
  GTECH_XOR2 U134 ( .A(n274), .B(n276), .Z(n271) );
  GTECH_AND_NOT U135 ( .A(n277), .B(n278), .Z(n274) );
  GTECH_XOR2 U136 ( .A(n279), .B(n280), .Z(sum[8]) );
  GTECH_MUX2 U137 ( .A(n281), .B(n282), .S(n283), .Z(sum[7]) );
  GTECH_XOR2 U138 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_AND_NOT U139 ( .A(n286), .B(n287), .Z(n285) );
  GTECH_OAI21 U140 ( .A(b[6]), .B(a[6]), .C(n288), .Z(n286) );
  GTECH_XOR2 U141 ( .A(n284), .B(n289), .Z(n281) );
  GTECH_XOR2 U142 ( .A(n290), .B(b[7]), .Z(n284) );
  GTECH_AO21 U143 ( .A(n291), .B(n287), .C(n292), .Z(sum[6]) );
  GTECH_NOT U144 ( .A(n293), .Z(n292) );
  GTECH_MUX2 U145 ( .A(n294), .B(n295), .S(b[6]), .Z(n293) );
  GTECH_OR_NOT U146 ( .A(n291), .B(n296), .Z(n295) );
  GTECH_XNOR2 U147 ( .A(a[6]), .B(n291), .Z(n294) );
  GTECH_AO21 U148 ( .A(n297), .B(n298), .C(n288), .Z(n291) );
  GTECH_NAND2 U149 ( .A(n299), .B(n300), .Z(n288) );
  GTECH_NAND3 U150 ( .A(b[4]), .B(n301), .C(a[4]), .Z(n299) );
  GTECH_MUX2 U151 ( .A(n302), .B(n303), .S(n304), .Z(sum[5]) );
  GTECH_AND2 U152 ( .A(n300), .B(n301), .Z(n304) );
  GTECH_OAI22 U153 ( .A(a[4]), .B(n298), .C(b[4]), .D(n305), .Z(n303) );
  GTECH_OR_NOT U154 ( .A(n305), .B(n306), .Z(n302) );
  GTECH_OAI21 U155 ( .A(a[4]), .B(n298), .C(b[4]), .Z(n306) );
  GTECH_AND2 U156 ( .A(a[4]), .B(n298), .Z(n305) );
  GTECH_XNOR2 U157 ( .A(n298), .B(n307), .Z(sum[4]) );
  GTECH_NOT U158 ( .A(n283), .Z(n298) );
  GTECH_MUX2 U159 ( .A(n308), .B(n309), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U160 ( .A(n310), .B(n311), .Z(n309) );
  GTECH_XNOR2 U161 ( .A(n312), .B(n310), .Z(n308) );
  GTECH_XNOR2 U162 ( .A(a[3]), .B(b[3]), .Z(n310) );
  GTECH_OA22 U163 ( .A(a[2]), .B(n313), .C(b[2]), .D(n314), .Z(n312) );
  GTECH_AND2 U164 ( .A(a[2]), .B(n313), .Z(n314) );
  GTECH_MUX2 U165 ( .A(n315), .B(n316), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U166 ( .A(n317), .B(n318), .Z(n316) );
  GTECH_XOR2 U167 ( .A(n317), .B(n313), .Z(n315) );
  GTECH_AO21 U168 ( .A(n319), .B(n320), .C(n321), .Z(n313) );
  GTECH_XOR2 U169 ( .A(a[2]), .B(b[2]), .Z(n317) );
  GTECH_MUX2 U170 ( .A(n322), .B(n323), .S(n324), .Z(sum[1]) );
  GTECH_AND_NOT U171 ( .A(n319), .B(n321), .Z(n324) );
  GTECH_OAI21 U172 ( .A(cin), .B(n320), .C(n325), .Z(n323) );
  GTECH_AO21 U173 ( .A(n325), .B(cin), .C(n320), .Z(n322) );
  GTECH_MUX2 U174 ( .A(n326), .B(n327), .S(n328), .Z(sum[15]) );
  GTECH_XOR2 U175 ( .A(n329), .B(n330), .Z(n327) );
  GTECH_XNOR2 U176 ( .A(n329), .B(n331), .Z(n326) );
  GTECH_AND_NOT U177 ( .A(n332), .B(n333), .Z(n331) );
  GTECH_OAI21 U178 ( .A(b[14]), .B(a[14]), .C(n334), .Z(n332) );
  GTECH_XOR2 U179 ( .A(a[15]), .B(b[15]), .Z(n329) );
  GTECH_AO21 U180 ( .A(n335), .B(n333), .C(n336), .Z(sum[14]) );
  GTECH_NOT U181 ( .A(n337), .Z(n336) );
  GTECH_MUX2 U182 ( .A(n338), .B(n339), .S(b[14]), .Z(n337) );
  GTECH_OR_NOT U183 ( .A(n335), .B(n340), .Z(n339) );
  GTECH_XNOR2 U184 ( .A(a[14]), .B(n335), .Z(n338) );
  GTECH_AO21 U185 ( .A(n341), .B(n328), .C(n334), .Z(n335) );
  GTECH_AO21 U186 ( .A(n342), .B(n343), .C(n344), .Z(n334) );
  GTECH_MUX2 U187 ( .A(n345), .B(n346), .S(n347), .Z(sum[13]) );
  GTECH_AND_NOT U188 ( .A(n342), .B(n344), .Z(n347) );
  GTECH_OAI21 U189 ( .A(a[12]), .B(n328), .C(n348), .Z(n346) );
  GTECH_AO21 U190 ( .A(n328), .B(a[12]), .C(b[12]), .Z(n348) );
  GTECH_AO21 U191 ( .A(n349), .B(n328), .C(n343), .Z(n345) );
  GTECH_XNOR2 U192 ( .A(n328), .B(n350), .Z(sum[12]) );
  GTECH_MUX2 U193 ( .A(n351), .B(n352), .S(n280), .Z(sum[11]) );
  GTECH_XOR2 U194 ( .A(n353), .B(n354), .Z(n352) );
  GTECH_XNOR2 U195 ( .A(n353), .B(n355), .Z(n351) );
  GTECH_AND_NOT U196 ( .A(n356), .B(n357), .Z(n355) );
  GTECH_OAI21 U197 ( .A(b[10]), .B(a[10]), .C(n358), .Z(n356) );
  GTECH_NOT U198 ( .A(n359), .Z(n358) );
  GTECH_OAI21 U199 ( .A(n275), .B(n278), .C(n277), .Z(n359) );
  GTECH_XOR2 U200 ( .A(a[11]), .B(b[11]), .Z(n353) );
  GTECH_AO21 U201 ( .A(n360), .B(n357), .C(n361), .Z(sum[10]) );
  GTECH_NOT U202 ( .A(n362), .Z(n361) );
  GTECH_MUX2 U203 ( .A(n363), .B(n364), .S(b[10]), .Z(n362) );
  GTECH_OR_NOT U204 ( .A(n360), .B(n365), .Z(n364) );
  GTECH_XNOR2 U205 ( .A(a[10]), .B(n360), .Z(n363) );
  GTECH_AO21 U206 ( .A(n366), .B(n280), .C(n367), .Z(n360) );
  GTECH_AO21 U207 ( .A(n275), .B(n277), .C(n278), .Z(n367) );
  GTECH_NOT U208 ( .A(n273), .Z(n280) );
  GTECH_XNOR2 U209 ( .A(cin), .B(n368), .Z(sum[0]) );
  GTECH_NOT U210 ( .A(n369), .Z(cout) );
  GTECH_MUX2 U211 ( .A(n350), .B(n370), .S(n328), .Z(n369) );
  GTECH_MUX2 U212 ( .A(n371), .B(n279), .S(n273), .Z(n328) );
  GTECH_MUX2 U213 ( .A(n372), .B(n307), .S(n283), .Z(n273) );
  GTECH_MUX2 U214 ( .A(n368), .B(n373), .S(cin), .Z(n283) );
  GTECH_AOI22 U215 ( .A(n311), .B(a[3]), .C(n374), .D(b[3]), .Z(n373) );
  GTECH_OR2 U216 ( .A(a[3]), .B(n311), .Z(n374) );
  GTECH_AO21 U217 ( .A(n318), .B(a[2]), .C(n375), .Z(n311) );
  GTECH_NOT U218 ( .A(n376), .Z(n375) );
  GTECH_OAI21 U219 ( .A(a[2]), .B(n318), .C(b[2]), .Z(n376) );
  GTECH_AO21 U220 ( .A(n325), .B(n319), .C(n321), .Z(n318) );
  GTECH_AND2 U221 ( .A(b[1]), .B(a[1]), .Z(n321) );
  GTECH_OR2 U222 ( .A(a[1]), .B(b[1]), .Z(n319) );
  GTECH_OR_NOT U223 ( .A(n320), .B(n325), .Z(n368) );
  GTECH_OR2 U224 ( .A(a[0]), .B(b[0]), .Z(n325) );
  GTECH_AND2 U225 ( .A(b[0]), .B(a[0]), .Z(n320) );
  GTECH_XNOR2 U226 ( .A(a[4]), .B(b[4]), .Z(n307) );
  GTECH_AOI2N2 U227 ( .A(n377), .B(b[7]), .C(n289), .D(n290), .Z(n372) );
  GTECH_NAND2 U228 ( .A(n290), .B(n289), .Z(n377) );
  GTECH_AND_NOT U229 ( .A(n378), .B(n287), .Z(n289) );
  GTECH_AND_NOT U230 ( .A(b[6]), .B(n296), .Z(n287) );
  GTECH_NOT U231 ( .A(a[6]), .Z(n296) );
  GTECH_OAI21 U232 ( .A(a[6]), .B(b[6]), .C(n297), .Z(n378) );
  GTECH_NAND2 U233 ( .A(n379), .B(n300), .Z(n297) );
  GTECH_NAND2 U234 ( .A(a[5]), .B(b[5]), .Z(n300) );
  GTECH_OAI21 U235 ( .A(a[4]), .B(b[4]), .C(n301), .Z(n379) );
  GTECH_OR2 U236 ( .A(b[5]), .B(a[5]), .Z(n301) );
  GTECH_NOT U237 ( .A(a[7]), .Z(n290) );
  GTECH_AND_NOT U238 ( .A(n276), .B(n275), .Z(n279) );
  GTECH_AND2 U239 ( .A(b[8]), .B(a[8]), .Z(n275) );
  GTECH_OA22 U240 ( .A(b[11]), .B(n380), .C(a[11]), .D(n354), .Z(n371) );
  GTECH_AND2 U241 ( .A(a[11]), .B(n354), .Z(n380) );
  GTECH_OR_NOT U242 ( .A(n357), .B(n381), .Z(n354) );
  GTECH_OAI21 U243 ( .A(a[10]), .B(b[10]), .C(n366), .Z(n381) );
  GTECH_AO21 U244 ( .A(n276), .B(n277), .C(n278), .Z(n366) );
  GTECH_AND2 U245 ( .A(a[9]), .B(b[9]), .Z(n278) );
  GTECH_OR2 U246 ( .A(b[9]), .B(a[9]), .Z(n277) );
  GTECH_OR2 U247 ( .A(a[8]), .B(b[8]), .Z(n276) );
  GTECH_AND_NOT U248 ( .A(b[10]), .B(n365), .Z(n357) );
  GTECH_NOT U249 ( .A(a[10]), .Z(n365) );
  GTECH_AOI21 U250 ( .A(n330), .B(a[15]), .C(n382), .Z(n370) );
  GTECH_NOT U251 ( .A(n383), .Z(n382) );
  GTECH_OAI21 U252 ( .A(a[15]), .B(n330), .C(b[15]), .Z(n383) );
  GTECH_OR_NOT U253 ( .A(n333), .B(n384), .Z(n330) );
  GTECH_OAI21 U254 ( .A(a[14]), .B(b[14]), .C(n341), .Z(n384) );
  GTECH_AO21 U255 ( .A(n342), .B(n349), .C(n344), .Z(n341) );
  GTECH_AND2 U256 ( .A(a[13]), .B(b[13]), .Z(n344) );
  GTECH_OR2 U257 ( .A(a[13]), .B(b[13]), .Z(n342) );
  GTECH_AND_NOT U258 ( .A(b[14]), .B(n340), .Z(n333) );
  GTECH_NOT U259 ( .A(a[14]), .Z(n340) );
  GTECH_OR_NOT U260 ( .A(n343), .B(n349), .Z(n350) );
  GTECH_OR2 U261 ( .A(b[12]), .B(a[12]), .Z(n349) );
  GTECH_AND2 U262 ( .A(a[12]), .B(b[12]), .Z(n343) );
endmodule

