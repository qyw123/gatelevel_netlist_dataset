
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142;

  GTECH_XOR2 U90 ( .A(n71), .B(n72), .Z(sum[9]) );
  GTECH_XOR2 U91 ( .A(n73), .B(n74), .Z(sum[8]) );
  GTECH_NOT U92 ( .A(n75), .Z(sum[7]) );
  GTECH_XOR2 U93 ( .A(n76), .B(n77), .Z(n75) );
  GTECH_AOI21 U94 ( .A(n78), .B(n79), .C(n80), .Z(n77) );
  GTECH_XOR2 U95 ( .A(n79), .B(n78), .Z(sum[6]) );
  GTECH_OAI2N2 U96 ( .A(n81), .B(n82), .C(n83), .D(n84), .Z(n78) );
  GTECH_XOR2 U97 ( .A(n84), .B(n83), .Z(sum[5]) );
  GTECH_OAI2N2 U98 ( .A(n85), .B(n86), .C(a[4]), .D(b[4]), .Z(n83) );
  GTECH_XOR2 U99 ( .A(n86), .B(n85), .Z(sum[4]) );
  GTECH_NOT U100 ( .A(n87), .Z(n86) );
  GTECH_XOR2 U101 ( .A(n88), .B(n89), .Z(sum[3]) );
  GTECH_AOI21 U102 ( .A(n90), .B(n91), .C(n92), .Z(n89) );
  GTECH_NOT U103 ( .A(n93), .Z(n88) );
  GTECH_XOR2 U104 ( .A(n91), .B(n90), .Z(sum[2]) );
  GTECH_AO21 U105 ( .A(n94), .B(n95), .C(n96), .Z(n90) );
  GTECH_XOR2 U106 ( .A(n95), .B(n94), .Z(sum[1]) );
  GTECH_NOT U107 ( .A(n97), .Z(n94) );
  GTECH_AOI22 U108 ( .A(n98), .B(cin), .C(a[0]), .D(b[0]), .Z(n97) );
  GTECH_XOR2 U109 ( .A(n99), .B(n100), .Z(sum[15]) );
  GTECH_AOI21 U110 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_XOR2 U111 ( .A(n102), .B(n101), .Z(sum[14]) );
  GTECH_OAI2N2 U112 ( .A(n104), .B(n105), .C(n106), .D(n107), .Z(n101) );
  GTECH_XOR2 U113 ( .A(n107), .B(n106), .Z(sum[13]) );
  GTECH_NOT U114 ( .A(n108), .Z(n106) );
  GTECH_AOI22 U115 ( .A(cout), .B(n109), .C(a[12]), .D(b[12]), .Z(n108) );
  GTECH_XOR2 U116 ( .A(n109), .B(cout), .Z(sum[12]) );
  GTECH_XOR2 U117 ( .A(n110), .B(n111), .Z(sum[11]) );
  GTECH_AOI21 U118 ( .A(n112), .B(n113), .C(n114), .Z(n111) );
  GTECH_XOR2 U119 ( .A(n113), .B(n112), .Z(sum[10]) );
  GTECH_OAI2N2 U120 ( .A(n115), .B(n116), .C(n72), .D(n71), .Z(n112) );
  GTECH_AO21 U121 ( .A(n74), .B(n73), .C(n117), .Z(n72) );
  GTECH_XOR2 U122 ( .A(cin), .B(n98), .Z(sum[0]) );
  GTECH_AO21 U123 ( .A(n74), .B(n118), .C(n119), .Z(cout) );
  GTECH_OAI21 U124 ( .A(n85), .B(n120), .C(n121), .Z(n74) );
  GTECH_AND2 U125 ( .A(n122), .B(n123), .Z(n85) );
  GTECH_NAND4 U126 ( .A(n124), .B(n98), .C(cin), .D(n125), .Z(n122) );
  GTECH_AND3 U127 ( .A(n91), .B(n95), .C(n93), .Z(n125) );
  GTECH_AND4 U128 ( .A(n126), .B(n124), .C(n118), .D(n127), .Z(Pm) );
  GTECH_AND4 U129 ( .A(n98), .B(n93), .C(n91), .D(n95), .Z(n127) );
  GTECH_XOR2 U130 ( .A(a[0]), .B(b[0]), .Z(n98) );
  GTECH_AO21 U131 ( .A(n128), .B(n118), .C(n119), .Z(Gm) );
  GTECH_OAI2N2 U132 ( .A(n129), .B(n99), .C(b[15]), .D(a[15]), .Z(n119) );
  GTECH_NOT U133 ( .A(n130), .Z(n99) );
  GTECH_AOI21 U134 ( .A(n131), .B(n102), .C(n103), .Z(n129) );
  GTECH_AND2 U135 ( .A(a[14]), .B(b[14]), .Z(n103) );
  GTECH_OAI21 U136 ( .A(n104), .B(n105), .C(n132), .Z(n131) );
  GTECH_NAND3 U137 ( .A(a[12]), .B(n107), .C(b[12]), .Z(n132) );
  GTECH_AND4 U138 ( .A(n109), .B(n130), .C(n102), .D(n107), .Z(n118) );
  GTECH_XOR2 U139 ( .A(n105), .B(n104), .Z(n107) );
  GTECH_NOT U140 ( .A(b[13]), .Z(n104) );
  GTECH_NOT U141 ( .A(a[13]), .Z(n105) );
  GTECH_XOR2 U142 ( .A(a[14]), .B(b[14]), .Z(n102) );
  GTECH_XOR2 U143 ( .A(a[15]), .B(b[15]), .Z(n130) );
  GTECH_XOR2 U144 ( .A(a[12]), .B(b[12]), .Z(n109) );
  GTECH_OAI21 U145 ( .A(n123), .B(n120), .C(n121), .Z(n128) );
  GTECH_AOI2N2 U146 ( .A(b[11]), .B(a[11]), .C(n133), .D(n110), .Z(n121) );
  GTECH_NOT U147 ( .A(n134), .Z(n110) );
  GTECH_AOI21 U148 ( .A(n135), .B(n113), .C(n114), .Z(n133) );
  GTECH_AND2 U149 ( .A(a[10]), .B(b[10]), .Z(n114) );
  GTECH_OAI2N2 U150 ( .A(n115), .B(n116), .C(n71), .D(n117), .Z(n135) );
  GTECH_AND2 U151 ( .A(a[8]), .B(b[8]), .Z(n117) );
  GTECH_NOT U152 ( .A(a[9]), .Z(n116) );
  GTECH_NOT U153 ( .A(b[9]), .Z(n115) );
  GTECH_NOT U154 ( .A(n126), .Z(n120) );
  GTECH_AND4 U155 ( .A(n73), .B(n134), .C(n113), .D(n71), .Z(n126) );
  GTECH_XOR2 U156 ( .A(a[9]), .B(b[9]), .Z(n71) );
  GTECH_XOR2 U157 ( .A(a[10]), .B(b[10]), .Z(n113) );
  GTECH_XOR2 U158 ( .A(a[11]), .B(b[11]), .Z(n134) );
  GTECH_XOR2 U159 ( .A(a[8]), .B(b[8]), .Z(n73) );
  GTECH_AOI222 U160 ( .A(n124), .B(n136), .C(b[7]), .D(a[7]), .E(n76), .F(n137), .Z(n123) );
  GTECH_AO21 U161 ( .A(n138), .B(n79), .C(n80), .Z(n137) );
  GTECH_AND2 U162 ( .A(a[6]), .B(b[6]), .Z(n80) );
  GTECH_OAI21 U163 ( .A(n81), .B(n82), .C(n139), .Z(n138) );
  GTECH_NAND3 U164 ( .A(a[4]), .B(n84), .C(b[4]), .Z(n139) );
  GTECH_NOT U165 ( .A(a[5]), .Z(n82) );
  GTECH_NOT U166 ( .A(b[5]), .Z(n81) );
  GTECH_AO21 U167 ( .A(b[3]), .B(a[3]), .C(n140), .Z(n136) );
  GTECH_OA21 U168 ( .A(n141), .B(n92), .C(n93), .Z(n140) );
  GTECH_XOR2 U169 ( .A(a[3]), .B(b[3]), .Z(n93) );
  GTECH_AND2 U170 ( .A(a[2]), .B(b[2]), .Z(n92) );
  GTECH_OA21 U171 ( .A(n142), .B(n96), .C(n91), .Z(n141) );
  GTECH_XOR2 U172 ( .A(a[2]), .B(b[2]), .Z(n91) );
  GTECH_AND2 U173 ( .A(a[1]), .B(b[1]), .Z(n96) );
  GTECH_AND3 U174 ( .A(a[0]), .B(n95), .C(b[0]), .Z(n142) );
  GTECH_XOR2 U175 ( .A(a[1]), .B(b[1]), .Z(n95) );
  GTECH_AND4 U176 ( .A(n87), .B(n84), .C(n79), .D(n76), .Z(n124) );
  GTECH_XOR2 U177 ( .A(a[7]), .B(b[7]), .Z(n76) );
  GTECH_XOR2 U178 ( .A(a[6]), .B(b[6]), .Z(n79) );
  GTECH_XOR2 U179 ( .A(a[5]), .B(b[5]), .Z(n84) );
  GTECH_XOR2 U180 ( .A(a[4]), .B(b[4]), .Z(n87) );
endmodule

