
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369;

  GTECH_MUX2 U132 ( .A(n271), .B(n272), .S(n273), .Z(sum[9]) );
  GTECH_XNOR2 U133 ( .A(n274), .B(n275), .Z(n272) );
  GTECH_XOR2 U134 ( .A(n274), .B(n276), .Z(n271) );
  GTECH_AND_NOT U135 ( .A(n277), .B(n278), .Z(n274) );
  GTECH_NAND2 U136 ( .A(n279), .B(n280), .Z(sum[8]) );
  GTECH_AO21 U137 ( .A(n275), .B(n276), .C(n273), .Z(n279) );
  GTECH_MUX2 U138 ( .A(n281), .B(n282), .S(n283), .Z(sum[7]) );
  GTECH_XNOR2 U139 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_XOR2 U140 ( .A(n284), .B(n286), .Z(n281) );
  GTECH_OA21 U141 ( .A(n287), .B(n288), .C(n289), .Z(n286) );
  GTECH_XNOR2 U142 ( .A(a[7]), .B(b[7]), .Z(n284) );
  GTECH_MUX2 U143 ( .A(n290), .B(n291), .S(n283), .Z(sum[6]) );
  GTECH_XNOR2 U144 ( .A(n292), .B(n293), .Z(n291) );
  GTECH_XNOR2 U145 ( .A(n288), .B(n292), .Z(n290) );
  GTECH_AND_NOT U146 ( .A(n289), .B(n287), .Z(n292) );
  GTECH_AOI21 U147 ( .A(n294), .B(n295), .C(n296), .Z(n288) );
  GTECH_MUX2 U148 ( .A(n297), .B(n298), .S(n299), .Z(sum[5]) );
  GTECH_AND_NOT U149 ( .A(n294), .B(n296), .Z(n299) );
  GTECH_OAI21 U150 ( .A(n295), .B(n283), .C(n300), .Z(n298) );
  GTECH_AO21 U151 ( .A(n300), .B(n283), .C(n295), .Z(n297) );
  GTECH_XOR2 U152 ( .A(n301), .B(n302), .Z(sum[4]) );
  GTECH_MUX2 U153 ( .A(n303), .B(n304), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U154 ( .A(n305), .B(n306), .Z(n304) );
  GTECH_XOR2 U155 ( .A(n305), .B(n307), .Z(n303) );
  GTECH_OA21 U156 ( .A(n308), .B(n309), .C(n310), .Z(n307) );
  GTECH_XNOR2 U157 ( .A(a[3]), .B(b[3]), .Z(n305) );
  GTECH_MUX2 U158 ( .A(n311), .B(n312), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U159 ( .A(n313), .B(n314), .Z(n312) );
  GTECH_XNOR2 U160 ( .A(n309), .B(n313), .Z(n311) );
  GTECH_AND_NOT U161 ( .A(n310), .B(n308), .Z(n313) );
  GTECH_AOI21 U162 ( .A(n315), .B(n316), .C(n317), .Z(n309) );
  GTECH_MUX2 U163 ( .A(n318), .B(n319), .S(n320), .Z(sum[1]) );
  GTECH_AND_NOT U164 ( .A(n315), .B(n317), .Z(n320) );
  GTECH_OAI21 U165 ( .A(cin), .B(n316), .C(n321), .Z(n319) );
  GTECH_AO21 U166 ( .A(n321), .B(cin), .C(n316), .Z(n318) );
  GTECH_AND_NOT U167 ( .A(b[0]), .B(n322), .Z(n316) );
  GTECH_MUX2 U168 ( .A(n323), .B(n324), .S(n325), .Z(sum[15]) );
  GTECH_XOR2 U169 ( .A(n326), .B(n327), .Z(n324) );
  GTECH_XOR2 U170 ( .A(n328), .B(n327), .Z(n323) );
  GTECH_XOR2 U171 ( .A(a[15]), .B(b[15]), .Z(n327) );
  GTECH_OA21 U172 ( .A(n329), .B(n330), .C(n331), .Z(n328) );
  GTECH_MUX2 U173 ( .A(n332), .B(n333), .S(n325), .Z(sum[14]) );
  GTECH_XNOR2 U174 ( .A(n334), .B(n335), .Z(n333) );
  GTECH_XNOR2 U175 ( .A(n334), .B(n330), .Z(n332) );
  GTECH_OA21 U176 ( .A(n336), .B(n337), .C(n338), .Z(n330) );
  GTECH_OAI21 U177 ( .A(a[14]), .B(b[14]), .C(n339), .Z(n334) );
  GTECH_NOT U178 ( .A(n329), .Z(n339) );
  GTECH_MUX2 U179 ( .A(n340), .B(n341), .S(n325), .Z(sum[13]) );
  GTECH_XOR2 U180 ( .A(n342), .B(n343), .Z(n341) );
  GTECH_XNOR2 U181 ( .A(n343), .B(n337), .Z(n340) );
  GTECH_OAI21 U182 ( .A(a[13]), .B(b[13]), .C(n344), .Z(n343) );
  GTECH_OR_NOT U183 ( .A(n345), .B(n346), .Z(sum[12]) );
  GTECH_OAI21 U184 ( .A(n337), .B(n342), .C(n325), .Z(n346) );
  GTECH_MUX2 U185 ( .A(n347), .B(n348), .S(n273), .Z(sum[11]) );
  GTECH_XOR2 U186 ( .A(n349), .B(n350), .Z(n348) );
  GTECH_OA21 U187 ( .A(n351), .B(n352), .C(n353), .Z(n350) );
  GTECH_NOR2 U188 ( .A(b[10]), .B(a[10]), .Z(n351) );
  GTECH_XNOR2 U189 ( .A(n349), .B(n354), .Z(n347) );
  GTECH_XNOR2 U190 ( .A(a[11]), .B(b[11]), .Z(n349) );
  GTECH_MUX2 U191 ( .A(n355), .B(n356), .S(n273), .Z(sum[10]) );
  GTECH_XOR2 U192 ( .A(n357), .B(n352), .Z(n356) );
  GTECH_AOI21 U193 ( .A(n277), .B(n358), .C(n278), .Z(n352) );
  GTECH_NOT U194 ( .A(n275), .Z(n358) );
  GTECH_XNOR2 U195 ( .A(n357), .B(n359), .Z(n355) );
  GTECH_OAI21 U196 ( .A(b[10]), .B(a[10]), .C(n353), .Z(n357) );
  GTECH_XNOR2 U197 ( .A(cin), .B(n360), .Z(sum[0]) );
  GTECH_AO21 U198 ( .A(n361), .B(n325), .C(n345), .Z(cout) );
  GTECH_NOR3 U199 ( .A(n337), .B(n342), .C(n325), .Z(n345) );
  GTECH_ADD_AB U200 ( .A(b[12]), .B(a[12]), .COUT(n337) );
  GTECH_OAI21 U201 ( .A(n362), .B(n273), .C(n280), .Z(n325) );
  GTECH_NAND3 U202 ( .A(n275), .B(n276), .C(n273), .Z(n280) );
  GTECH_NAND2 U203 ( .A(b[8]), .B(a[8]), .Z(n275) );
  GTECH_MUX2 U204 ( .A(n301), .B(n363), .S(n283), .Z(n273) );
  GTECH_NOT U205 ( .A(n302), .Z(n283) );
  GTECH_MUX2 U206 ( .A(n360), .B(n364), .S(cin), .Z(n302) );
  GTECH_AOI21 U207 ( .A(n306), .B(a[3]), .C(n365), .Z(n364) );
  GTECH_OA21 U208 ( .A(a[3]), .B(n306), .C(b[3]), .Z(n365) );
  GTECH_OAI21 U209 ( .A(n314), .B(n308), .C(n310), .Z(n306) );
  GTECH_NAND2 U210 ( .A(b[2]), .B(a[2]), .Z(n310) );
  GTECH_NOR2 U211 ( .A(a[2]), .B(b[2]), .Z(n308) );
  GTECH_AOI21 U212 ( .A(n321), .B(n315), .C(n317), .Z(n314) );
  GTECH_ADD_AB U213 ( .A(a[1]), .B(b[1]), .COUT(n317) );
  GTECH_OR2 U214 ( .A(b[1]), .B(a[1]), .Z(n315) );
  GTECH_OR_NOT U215 ( .A(b[0]), .B(n322), .Z(n321) );
  GTECH_NOT U216 ( .A(a[0]), .Z(n322) );
  GTECH_XNOR2 U217 ( .A(a[0]), .B(b[0]), .Z(n360) );
  GTECH_AOI21 U218 ( .A(n285), .B(a[7]), .C(n366), .Z(n363) );
  GTECH_OA21 U219 ( .A(a[7]), .B(n285), .C(b[7]), .Z(n366) );
  GTECH_OAI21 U220 ( .A(n293), .B(n287), .C(n289), .Z(n285) );
  GTECH_NAND2 U221 ( .A(b[6]), .B(a[6]), .Z(n289) );
  GTECH_NOR2 U222 ( .A(a[6]), .B(b[6]), .Z(n287) );
  GTECH_AOI21 U223 ( .A(n300), .B(n294), .C(n296), .Z(n293) );
  GTECH_ADD_AB U224 ( .A(b[5]), .B(a[5]), .COUT(n296) );
  GTECH_OR2 U225 ( .A(a[5]), .B(b[5]), .Z(n294) );
  GTECH_OR_NOT U226 ( .A(n295), .B(n300), .Z(n301) );
  GTECH_OR2 U227 ( .A(b[4]), .B(a[4]), .Z(n300) );
  GTECH_ADD_AB U228 ( .A(b[4]), .B(a[4]), .COUT(n295) );
  GTECH_AOI21 U229 ( .A(n354), .B(a[11]), .C(n367), .Z(n362) );
  GTECH_OA21 U230 ( .A(a[11]), .B(n354), .C(b[11]), .Z(n367) );
  GTECH_NAND2 U231 ( .A(n368), .B(n353), .Z(n354) );
  GTECH_NAND2 U232 ( .A(b[10]), .B(a[10]), .Z(n353) );
  GTECH_OAI21 U233 ( .A(a[10]), .B(b[10]), .C(n359), .Z(n368) );
  GTECH_AO21 U234 ( .A(n276), .B(n277), .C(n278), .Z(n359) );
  GTECH_ADD_AB U235 ( .A(b[9]), .B(a[9]), .COUT(n278) );
  GTECH_OR2 U236 ( .A(a[9]), .B(b[9]), .Z(n277) );
  GTECH_OR2 U237 ( .A(a[8]), .B(b[8]), .Z(n276) );
  GTECH_ADD_ABC U238 ( .A(a[15]), .B(n326), .C(b[15]), .COUT(n361) );
  GTECH_OA21 U239 ( .A(n329), .B(n335), .C(n331), .Z(n326) );
  GTECH_OR2 U240 ( .A(b[14]), .B(a[14]), .Z(n331) );
  GTECH_AOI21 U241 ( .A(n344), .B(n342), .C(n369), .Z(n335) );
  GTECH_NOT U242 ( .A(n338), .Z(n369) );
  GTECH_OR2 U243 ( .A(b[13]), .B(a[13]), .Z(n338) );
  GTECH_NOR2 U244 ( .A(a[12]), .B(b[12]), .Z(n342) );
  GTECH_NOT U245 ( .A(n336), .Z(n344) );
  GTECH_ADD_AB U246 ( .A(a[13]), .B(b[13]), .COUT(n336) );
  GTECH_ADD_AB U247 ( .A(a[14]), .B(b[14]), .COUT(n329) );
endmodule

