
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134;

  GTECH_XOR2 U87 ( .A(n68), .B(n69), .Z(sum[9]) );
  GTECH_XOR2 U88 ( .A(n70), .B(n71), .Z(sum[8]) );
  GTECH_XOR2 U89 ( .A(n72), .B(n73), .Z(sum[7]) );
  GTECH_AOI21 U90 ( .A(n74), .B(n75), .C(n76), .Z(n73) );
  GTECH_NOT U91 ( .A(n77), .Z(n72) );
  GTECH_XOR2 U92 ( .A(n75), .B(n74), .Z(sum[6]) );
  GTECH_AO22 U93 ( .A(n78), .B(n79), .C(b[5]), .D(a[5]), .Z(n74) );
  GTECH_XOR2 U94 ( .A(n79), .B(n78), .Z(sum[5]) );
  GTECH_AO22 U95 ( .A(n80), .B(n81), .C(b[4]), .D(a[4]), .Z(n78) );
  GTECH_XOR2 U96 ( .A(n81), .B(n80), .Z(sum[4]) );
  GTECH_XOR2 U97 ( .A(n82), .B(n83), .Z(sum[3]) );
  GTECH_AOI21 U98 ( .A(n84), .B(n85), .C(n86), .Z(n83) );
  GTECH_XOR2 U99 ( .A(n85), .B(n84), .Z(sum[2]) );
  GTECH_OAI2N2 U100 ( .A(n87), .B(n88), .C(b[1]), .D(a[1]), .Z(n84) );
  GTECH_XOR2 U101 ( .A(n88), .B(n87), .Z(sum[1]) );
  GTECH_AOI22 U102 ( .A(n89), .B(cin), .C(a[0]), .D(b[0]), .Z(n87) );
  GTECH_NOT U103 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U104 ( .A(n91), .B(n92), .Z(sum[15]) );
  GTECH_OA21 U105 ( .A(n93), .B(n94), .C(n95), .Z(n92) );
  GTECH_XOR2 U106 ( .A(n94), .B(n93), .Z(sum[14]) );
  GTECH_AOI22 U107 ( .A(b[13]), .B(a[13]), .C(n96), .D(n97), .Z(n93) );
  GTECH_XOR2 U108 ( .A(n97), .B(n96), .Z(sum[13]) );
  GTECH_AO22 U109 ( .A(a[12]), .B(b[12]), .C(cout), .D(n98), .Z(n96) );
  GTECH_XOR2 U110 ( .A(n98), .B(cout), .Z(sum[12]) );
  GTECH_XOR2 U111 ( .A(n99), .B(n100), .Z(sum[11]) );
  GTECH_OA21 U112 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_NOT U113 ( .A(n104), .Z(n99) );
  GTECH_XOR2 U114 ( .A(n102), .B(n101), .Z(sum[10]) );
  GTECH_OA21 U115 ( .A(n68), .B(n69), .C(n105), .Z(n101) );
  GTECH_AOI21 U116 ( .A(n70), .B(n71), .C(n106), .Z(n69) );
  GTECH_NOT U117 ( .A(n107), .Z(n68) );
  GTECH_NOT U118 ( .A(n108), .Z(n102) );
  GTECH_XOR2 U119 ( .A(cin), .B(n89), .Z(sum[0]) );
  GTECH_AO21 U120 ( .A(n109), .B(n71), .C(n110), .Z(cout) );
  GTECH_AO21 U121 ( .A(n111), .B(n80), .C(n112), .Z(n71) );
  GTECH_AO21 U122 ( .A(cin), .B(n113), .C(n114), .Z(n80) );
  GTECH_AND3 U123 ( .A(n111), .B(n113), .C(n109), .Z(Pm) );
  GTECH_AND5 U124 ( .A(n85), .B(n90), .C(n115), .D(n116), .E(n89), .Z(n113) );
  GTECH_XOR2 U125 ( .A(a[0]), .B(b[0]), .Z(n89) );
  GTECH_AO21 U126 ( .A(n109), .B(n117), .C(n110), .Z(Gm) );
  GTECH_OAI2N2 U127 ( .A(n118), .B(n91), .C(b[15]), .D(a[15]), .Z(n110) );
  GTECH_NOT U128 ( .A(n119), .Z(n91) );
  GTECH_OA21 U129 ( .A(n120), .B(n94), .C(n95), .Z(n118) );
  GTECH_NAND2 U130 ( .A(b[14]), .B(a[14]), .Z(n95) );
  GTECH_NOT U131 ( .A(n121), .Z(n94) );
  GTECH_AOI21 U132 ( .A(b[13]), .B(a[13]), .C(n122), .Z(n120) );
  GTECH_AND3 U133 ( .A(a[12]), .B(n97), .C(b[12]), .Z(n122) );
  GTECH_AO21 U134 ( .A(n111), .B(n114), .C(n112), .Z(n117) );
  GTECH_AO22 U135 ( .A(b[11]), .B(a[11]), .C(n123), .D(n104), .Z(n112) );
  GTECH_AO21 U136 ( .A(n124), .B(n108), .C(n125), .Z(n123) );
  GTECH_AO21 U137 ( .A(n106), .B(n107), .C(n126), .Z(n124) );
  GTECH_NOT U138 ( .A(n105), .Z(n126) );
  GTECH_AND2 U139 ( .A(b[8]), .B(a[8]), .Z(n106) );
  GTECH_NOT U140 ( .A(n127), .Z(n114) );
  GTECH_AOI222 U141 ( .A(a[7]), .B(b[7]), .C(n116), .D(n128), .E(n77), .F(n129), .Z(n127) );
  GTECH_AO21 U142 ( .A(n75), .B(n130), .C(n76), .Z(n129) );
  GTECH_AND2 U143 ( .A(b[6]), .B(a[6]), .Z(n76) );
  GTECH_AO22 U144 ( .A(a[4]), .B(n131), .C(b[5]), .D(a[5]), .Z(n130) );
  GTECH_AND2 U145 ( .A(n79), .B(b[4]), .Z(n131) );
  GTECH_OAI2N2 U146 ( .A(n132), .B(n82), .C(b[3]), .D(a[3]), .Z(n128) );
  GTECH_NOT U147 ( .A(n115), .Z(n82) );
  GTECH_XOR2 U148 ( .A(a[3]), .B(b[3]), .Z(n115) );
  GTECH_AOI21 U149 ( .A(n133), .B(n85), .C(n86), .Z(n132) );
  GTECH_AND2 U150 ( .A(b[2]), .B(a[2]), .Z(n86) );
  GTECH_XOR2 U151 ( .A(a[2]), .B(b[2]), .Z(n85) );
  GTECH_AO21 U152 ( .A(b[1]), .B(a[1]), .C(n134), .Z(n133) );
  GTECH_AND3 U153 ( .A(a[0]), .B(n90), .C(b[0]), .Z(n134) );
  GTECH_XOR2 U154 ( .A(a[1]), .B(b[1]), .Z(n90) );
  GTECH_AND4 U155 ( .A(n81), .B(n79), .C(n75), .D(n77), .Z(n116) );
  GTECH_XOR2 U156 ( .A(a[7]), .B(b[7]), .Z(n77) );
  GTECH_XOR2 U157 ( .A(a[6]), .B(b[6]), .Z(n75) );
  GTECH_XOR2 U158 ( .A(a[5]), .B(b[5]), .Z(n79) );
  GTECH_XOR2 U159 ( .A(a[4]), .B(b[4]), .Z(n81) );
  GTECH_AND4 U160 ( .A(n108), .B(n107), .C(n70), .D(n104), .Z(n111) );
  GTECH_XOR2 U161 ( .A(a[11]), .B(b[11]), .Z(n104) );
  GTECH_XOR2 U162 ( .A(a[8]), .B(b[8]), .Z(n70) );
  GTECH_OA21 U163 ( .A(a[9]), .B(b[9]), .C(n105), .Z(n107) );
  GTECH_NAND2 U164 ( .A(b[9]), .B(a[9]), .Z(n105) );
  GTECH_OA21 U165 ( .A(a[10]), .B(b[10]), .C(n103), .Z(n108) );
  GTECH_NOT U166 ( .A(n125), .Z(n103) );
  GTECH_AND2 U167 ( .A(b[10]), .B(a[10]), .Z(n125) );
  GTECH_AND4 U168 ( .A(n98), .B(n119), .C(n121), .D(n97), .Z(n109) );
  GTECH_XOR2 U169 ( .A(a[13]), .B(b[13]), .Z(n97) );
  GTECH_XOR2 U170 ( .A(a[14]), .B(b[14]), .Z(n121) );
  GTECH_XOR2 U171 ( .A(a[15]), .B(b[15]), .Z(n119) );
  GTECH_XOR2 U172 ( .A(a[12]), .B(b[12]), .Z(n98) );
endmodule

