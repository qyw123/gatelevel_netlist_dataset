
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n113, n114, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK2S Cntr_reg_0_ ( .J(n114), .K(n114), .TI(N14), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[0]), .QN(n338) );
  GTECH_FJK2S Cntr_reg_1_ ( .J(n114), .K(n114), .TI(N15), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK2S Cntr_reg_2_ ( .J(n114), .K(n114), .TI(N16), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK2S Cntr_reg_3_ ( .J(n114), .K(n114), .TI(N17), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK2S Cntr_reg_4_ ( .J(n114), .K(n114), .TI(N19), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK2S A_reg_16_ ( .J(n114), .K(n114), .TI(N42), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[16]), .QN(n355) );
  GTECH_FJK2S A_reg_15_ ( .J(n114), .K(n114), .TI(N42), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[15]), .QN(n354) );
  GTECH_FJK2S A_reg_14_ ( .J(n114), .K(n114), .TI(N39), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[14]), .QN(n353) );
  GTECH_FJK2S A_reg_13_ ( .J(n114), .K(n114), .TI(N38), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[13]), .QN(n352) );
  GTECH_FJK2S A_reg_12_ ( .J(n114), .K(n114), .TI(N37), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[12]), .QN(n351) );
  GTECH_FJK2S A_reg_11_ ( .J(n114), .K(n114), .TI(N36), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[11]), .QN(n350) );
  GTECH_FJK2S A_reg_10_ ( .J(n114), .K(n114), .TI(N35), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[10]), .QN(n349) );
  GTECH_FJK2S A_reg_9_ ( .J(n114), .K(n114), .TI(N34), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[9]), .QN(n348) );
  GTECH_FJK2S A_reg_8_ ( .J(n114), .K(n114), .TI(N33), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[8]), .QN(n347) );
  GTECH_FJK2S A_reg_7_ ( .J(n114), .K(n114), .TI(N32), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[7]), .QN(n346) );
  GTECH_FJK2S A_reg_6_ ( .J(n114), .K(n114), .TI(N31), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[6]), .QN(n345) );
  GTECH_FJK2S A_reg_5_ ( .J(n114), .K(n114), .TI(N30), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[5]), .QN(n344) );
  GTECH_FJK2S A_reg_4_ ( .J(n114), .K(n114), .TI(N29), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[4]), .QN(n343) );
  GTECH_FJK2S A_reg_3_ ( .J(n114), .K(n114), .TI(N28), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[3]), .QN(n342) );
  GTECH_FJK2S A_reg_2_ ( .J(n114), .K(n114), .TI(N27), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[2]), .QN(n341) );
  GTECH_FJK2S A_reg_1_ ( .J(n114), .K(n114), .TI(N26), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[1]), .QN(n340) );
  GTECH_FJK2S A_reg_0_ ( .J(n114), .K(n114), .TI(N25), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[0]), .QN(n339) );
  GTECH_FJK2S Prod_reg_0_ ( .J(n114), .K(n114), .TI(N82), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[0]), .QN(n10) );
  GTECH_FJK2S Prod_reg_18_ ( .J(n114), .K(n114), .TI(N100), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK2S Prod_reg_17_ ( .J(n114), .K(n114), .TI(N99), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[17]), .QN(n12) );
  GTECH_FJK2S Prod_reg_16_ ( .J(n114), .K(n114), .TI(N98), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[16]), .QN(n13) );
  GTECH_FJK2S Prod_reg_15_ ( .J(n114), .K(n114), .TI(N97), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[15]), .QN(n14) );
  GTECH_FJK2S Prod_reg_14_ ( .J(n114), .K(n114), .TI(N96), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[14]), .QN(n15) );
  GTECH_FJK2S Prod_reg_13_ ( .J(n114), .K(n114), .TI(N95), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[13]), .QN(n16) );
  GTECH_FJK2S Prod_reg_12_ ( .J(n114), .K(n114), .TI(N94), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[12]), .QN(n17) );
  GTECH_FJK2S Prod_reg_11_ ( .J(n114), .K(n114), .TI(N93), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[11]), .QN(n18) );
  GTECH_FJK2S Prod_reg_10_ ( .J(n114), .K(n114), .TI(N92), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[10]), .QN(n19) );
  GTECH_FJK2S Prod_reg_9_ ( .J(n114), .K(n114), .TI(N91), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[9]), .QN(n20) );
  GTECH_FJK2S Prod_reg_8_ ( .J(n114), .K(n114), .TI(N90), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[8]), .QN(n21) );
  GTECH_FJK2S Prod_reg_7_ ( .J(n114), .K(n114), .TI(N89), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[7]), .QN(n22) );
  GTECH_FJK2S Prod_reg_6_ ( .J(n114), .K(n114), .TI(N88), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[6]), .QN(n23) );
  GTECH_FJK2S Prod_reg_5_ ( .J(n114), .K(n114), .TI(N87), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[5]), .QN(n24) );
  GTECH_FJK2S Prod_reg_4_ ( .J(n114), .K(n114), .TI(N86), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[4]), .QN(n25) );
  GTECH_FJK2S Prod_reg_3_ ( .J(n114), .K(n114), .TI(N85), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[3]), .QN(n26) );
  GTECH_FJK2S Prod_reg_2_ ( .J(n114), .K(n114), .TI(N84), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[2]), .QN(n27) );
  GTECH_FJK2S Prod_reg_1_ ( .J(n114), .K(n114), .TI(N83), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[1]), .QN(n28) );
  GTECH_FJK2S Prod_reg_19_ ( .J(n114), .K(n114), .TI(N101), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK2S Prod_reg_33_ ( .J(n114), .K(n114), .TI(N116), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK2S Prod_reg_32_ ( .J(n114), .K(n114), .TI(N116), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK2S Prod_reg_31_ ( .J(n114), .K(n114), .TI(N113), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK2S Prod_reg_30_ ( .J(n114), .K(n114), .TI(N112), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK2S Prod_reg_29_ ( .J(n114), .K(n114), .TI(N111), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK2S Prod_reg_28_ ( .J(n114), .K(n114), .TI(N110), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK2S Prod_reg_27_ ( .J(n114), .K(n114), .TI(N109), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK2S Prod_reg_26_ ( .J(n114), .K(n114), .TI(N108), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK2S Prod_reg_25_ ( .J(n114), .K(n114), .TI(N107), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK2S Prod_reg_24_ ( .J(n114), .K(n114), .TI(N106), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK2S Prod_reg_23_ ( .J(n114), .K(n114), .TI(N105), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK2S Prod_reg_22_ ( .J(n114), .K(n114), .TI(N104), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK2S Prod_reg_21_ ( .J(n114), .K(n114), .TI(N103), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK2S Prod_reg_20_ ( .J(n114), .K(n114), .TI(N102), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK2S P_reg_31_ ( .J(n114), .K(n114), .TI(N152), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[31]) );
  GTECH_FJK2S P_reg_30_ ( .J(n114), .K(n114), .TI(N150), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[30]) );
  GTECH_FJK2S P_reg_29_ ( .J(n114), .K(n114), .TI(N149), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[29]) );
  GTECH_FJK2S P_reg_28_ ( .J(n114), .K(n114), .TI(N148), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[28]) );
  GTECH_FJK2S P_reg_27_ ( .J(n114), .K(n114), .TI(N147), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[27]) );
  GTECH_FJK2S P_reg_26_ ( .J(n114), .K(n114), .TI(N146), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[26]) );
  GTECH_FJK2S P_reg_25_ ( .J(n114), .K(n114), .TI(N145), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[25]) );
  GTECH_FJK2S P_reg_24_ ( .J(n114), .K(n114), .TI(N144), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[24]) );
  GTECH_FJK2S P_reg_23_ ( .J(n114), .K(n114), .TI(N143), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[23]) );
  GTECH_FJK2S P_reg_22_ ( .J(n114), .K(n114), .TI(N142), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[22]) );
  GTECH_FJK2S P_reg_21_ ( .J(n114), .K(n114), .TI(N141), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[21]) );
  GTECH_FJK2S P_reg_20_ ( .J(n114), .K(n114), .TI(N140), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[20]) );
  GTECH_FJK2S P_reg_19_ ( .J(n114), .K(n114), .TI(N139), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[19]) );
  GTECH_FJK2S P_reg_18_ ( .J(n114), .K(n114), .TI(N138), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[18]) );
  GTECH_FJK2S P_reg_17_ ( .J(n114), .K(n114), .TI(N137), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[17]) );
  GTECH_FJK2S P_reg_16_ ( .J(n114), .K(n114), .TI(N136), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[16]) );
  GTECH_FJK2S P_reg_15_ ( .J(n114), .K(n114), .TI(N135), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[15]) );
  GTECH_FJK2S P_reg_14_ ( .J(n114), .K(n114), .TI(N134), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[14]) );
  GTECH_FJK2S P_reg_13_ ( .J(n114), .K(n114), .TI(N133), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[13]) );
  GTECH_FJK2S P_reg_12_ ( .J(n114), .K(n114), .TI(N132), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[12]) );
  GTECH_FJK2S P_reg_11_ ( .J(n114), .K(n114), .TI(N131), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[11]) );
  GTECH_FJK2S P_reg_10_ ( .J(n114), .K(n114), .TI(N130), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[10]) );
  GTECH_FJK2S P_reg_9_ ( .J(n114), .K(n114), .TI(N129), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[9]) );
  GTECH_FJK2S P_reg_8_ ( .J(n114), .K(n114), .TI(N128), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[8]) );
  GTECH_FJK2S P_reg_7_ ( .J(n114), .K(n114), .TI(N127), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[7]) );
  GTECH_FJK2S P_reg_6_ ( .J(n114), .K(n114), .TI(N126), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[6]) );
  GTECH_FJK2S P_reg_5_ ( .J(n114), .K(n114), .TI(N125), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[5]) );
  GTECH_FJK2S P_reg_4_ ( .J(n114), .K(n114), .TI(N124), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[4]) );
  GTECH_FJK2S P_reg_3_ ( .J(n114), .K(n114), .TI(N123), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[3]) );
  GTECH_FJK2S P_reg_2_ ( .J(n114), .K(n114), .TI(N122), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[2]) );
  GTECH_FJK2S P_reg_1_ ( .J(n114), .K(n114), .TI(N121), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[1]) );
  GTECH_FJK2S P_reg_0_ ( .J(n114), .K(n114), .TI(N120), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U340 ( .Z(n114) );
  GTECH_ONE U341 ( .Z(n113) );
  GTECH_NOT U342 ( .A(n356), .Z(N99) );
  GTECH_AOI222 U343 ( .A(n357), .B(n358), .C(n359), .D(n360), .E(n361), .F(
        n362), .Z(n356) );
  GTECH_NOT U344 ( .A(n363), .Z(N98) );
  GTECH_AOI222 U345 ( .A(n359), .B(n364), .C(n365), .D(n366), .E(R[15]), .F(
        n367), .Z(n363) );
  GTECH_NAND2 U346 ( .A(n368), .B(n369), .Z(n365) );
  GTECH_OAI2N2 U347 ( .A(n13), .B(n370), .C(R[14]), .D(n367), .Z(N97) );
  GTECH_OAI2N2 U348 ( .A(n14), .B(n370), .C(R[13]), .D(n367), .Z(N96) );
  GTECH_OAI2N2 U349 ( .A(n15), .B(n370), .C(R[12]), .D(n367), .Z(N95) );
  GTECH_OAI2N2 U350 ( .A(n16), .B(n370), .C(R[11]), .D(n367), .Z(N94) );
  GTECH_OAI2N2 U351 ( .A(n17), .B(n370), .C(R[10]), .D(n367), .Z(N93) );
  GTECH_OAI2N2 U352 ( .A(n18), .B(n370), .C(R[9]), .D(n367), .Z(N92) );
  GTECH_OAI2N2 U353 ( .A(n19), .B(n370), .C(R[8]), .D(n367), .Z(N91) );
  GTECH_OAI2N2 U354 ( .A(n20), .B(n370), .C(R[7]), .D(n367), .Z(N90) );
  GTECH_OAI2N2 U355 ( .A(n21), .B(n370), .C(R[6]), .D(n367), .Z(N89) );
  GTECH_OAI2N2 U356 ( .A(n22), .B(n370), .C(R[5]), .D(n367), .Z(N88) );
  GTECH_OAI2N2 U357 ( .A(n23), .B(n370), .C(R[4]), .D(n367), .Z(N87) );
  GTECH_OAI2N2 U358 ( .A(n24), .B(n370), .C(R[3]), .D(n367), .Z(N86) );
  GTECH_OAI2N2 U359 ( .A(n25), .B(n370), .C(R[2]), .D(n367), .Z(N85) );
  GTECH_OAI2N2 U360 ( .A(n26), .B(n370), .C(R[1]), .D(n367), .Z(N84) );
  GTECH_OAI2N2 U361 ( .A(n27), .B(n370), .C(R[0]), .D(n367), .Z(N83) );
  GTECH_AND2 U362 ( .A(M[15]), .B(n367), .Z(N42) );
  GTECH_AND2 U363 ( .A(M[14]), .B(n367), .Z(N39) );
  GTECH_AND2 U364 ( .A(M[13]), .B(n367), .Z(N38) );
  GTECH_AND2 U365 ( .A(M[12]), .B(n367), .Z(N37) );
  GTECH_AND2 U366 ( .A(M[11]), .B(n367), .Z(N36) );
  GTECH_AND2 U367 ( .A(M[10]), .B(n367), .Z(N35) );
  GTECH_AND2 U368 ( .A(M[9]), .B(n367), .Z(N34) );
  GTECH_AND2 U369 ( .A(M[8]), .B(n367), .Z(N33) );
  GTECH_AND2 U370 ( .A(M[7]), .B(n367), .Z(N32) );
  GTECH_AND2 U371 ( .A(M[6]), .B(n367), .Z(N31) );
  GTECH_AND2 U372 ( .A(M[5]), .B(n367), .Z(N30) );
  GTECH_AND2 U373 ( .A(M[4]), .B(n367), .Z(N29) );
  GTECH_AND2 U374 ( .A(M[3]), .B(n367), .Z(N28) );
  GTECH_AND2 U375 ( .A(M[2]), .B(n367), .Z(N27) );
  GTECH_AND2 U376 ( .A(M[1]), .B(n367), .Z(N26) );
  GTECH_AND2 U377 ( .A(M[0]), .B(n367), .Z(N25) );
  GTECH_NOT U378 ( .A(n371), .Z(n367) );
  GTECH_NAND2 U379 ( .A(n371), .B(n372), .Z(N19) );
  GTECH_NAND3 U380 ( .A(n373), .B(n374), .C(n375), .Z(n372) );
  GTECH_NAND3 U381 ( .A(n376), .B(n377), .C(n370), .Z(N18) );
  GTECH_AND2 U382 ( .A(n375), .B(n378), .Z(N17) );
  GTECH_OAI21 U383 ( .A(n8), .B(n379), .C(n373), .Z(n378) );
  GTECH_AND2 U384 ( .A(n375), .B(n380), .Z(N16) );
  GTECH_OAI21 U385 ( .A(n7), .B(n381), .C(n382), .Z(n380) );
  GTECH_NOT U386 ( .A(n383), .Z(N152) );
  GTECH_AOI222 U387 ( .A(n384), .B(n385), .C(n386), .D(n387), .E(n388), .F(
        n389), .Z(n383) );
  GTECH_NAND2 U388 ( .A(n377), .B(n390), .Z(N151) );
  GTECH_NOT U389 ( .A(n391), .Z(N150) );
  GTECH_AOI222 U390 ( .A(n392), .B(n384), .C(n386), .D(n393), .E(n388), .F(
        n394), .Z(n391) );
  GTECH_MUX2 U391 ( .A(n395), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND2 U392 ( .A(n375), .B(n396), .Z(n395) );
  GTECH_NOT U393 ( .A(n397), .Z(N149) );
  GTECH_AOI222 U394 ( .A(n398), .B(n384), .C(n386), .D(n399), .E(n388), .F(
        n400), .Z(n397) );
  GTECH_NOT U395 ( .A(n401), .Z(N148) );
  GTECH_AOI222 U396 ( .A(n402), .B(n384), .C(n386), .D(n403), .E(n388), .F(
        n404), .Z(n401) );
  GTECH_NOT U397 ( .A(n405), .Z(N147) );
  GTECH_AOI222 U398 ( .A(n406), .B(n384), .C(n386), .D(n407), .E(n388), .F(
        n408), .Z(n405) );
  GTECH_NOT U399 ( .A(n409), .Z(N146) );
  GTECH_AOI222 U400 ( .A(n410), .B(n384), .C(n386), .D(n411), .E(n388), .F(
        n412), .Z(n409) );
  GTECH_NOT U401 ( .A(n413), .Z(N145) );
  GTECH_AOI222 U402 ( .A(n414), .B(n384), .C(n386), .D(n415), .E(n388), .F(
        n416), .Z(n413) );
  GTECH_NOT U403 ( .A(n417), .Z(N144) );
  GTECH_AOI222 U404 ( .A(n418), .B(n384), .C(n386), .D(n419), .E(n388), .F(
        n420), .Z(n417) );
  GTECH_NOT U405 ( .A(n421), .Z(N143) );
  GTECH_AOI222 U406 ( .A(n422), .B(n384), .C(n386), .D(n423), .E(n388), .F(
        n424), .Z(n421) );
  GTECH_NOT U407 ( .A(n425), .Z(N142) );
  GTECH_AOI222 U408 ( .A(n426), .B(n384), .C(n386), .D(n427), .E(n388), .F(
        n428), .Z(n425) );
  GTECH_NOT U409 ( .A(n429), .Z(N141) );
  GTECH_AOI222 U410 ( .A(n430), .B(n384), .C(n386), .D(n431), .E(n388), .F(
        n432), .Z(n429) );
  GTECH_NOT U411 ( .A(n433), .Z(N140) );
  GTECH_AOI222 U412 ( .A(n434), .B(n384), .C(n386), .D(n435), .E(n388), .F(
        n436), .Z(n433) );
  GTECH_NOT U413 ( .A(n437), .Z(N14) );
  GTECH_NAND2 U414 ( .A(n375), .B(n338), .Z(n437) );
  GTECH_NOT U415 ( .A(n438), .Z(N139) );
  GTECH_AOI222 U416 ( .A(n439), .B(n384), .C(n386), .D(n440), .E(n388), .F(
        n441), .Z(n438) );
  GTECH_NOT U417 ( .A(n442), .Z(N138) );
  GTECH_AOI222 U418 ( .A(n443), .B(n384), .C(n386), .D(n444), .E(n388), .F(
        n445), .Z(n442) );
  GTECH_NOT U419 ( .A(n446), .Z(N137) );
  GTECH_AOI222 U420 ( .A(n447), .B(n384), .C(n386), .D(n448), .E(n388), .F(
        n449), .Z(n446) );
  GTECH_NOT U421 ( .A(n450), .Z(N136) );
  GTECH_AOI222 U422 ( .A(n384), .B(n358), .C(n386), .D(n360), .E(n388), .F(
        n362), .Z(n450) );
  GTECH_NOT U423 ( .A(n451), .Z(n362) );
  GTECH_XNOR2 U424 ( .A(n452), .B(n453), .Z(n451) );
  GTECH_NOT U425 ( .A(n454), .Z(n452) );
  GTECH_NOT U426 ( .A(n455), .Z(n386) );
  GTECH_NOT U427 ( .A(n456), .Z(n358) );
  GTECH_XNOR2 U428 ( .A(n457), .B(n453), .Z(n456) );
  GTECH_NOT U429 ( .A(n458), .Z(n453) );
  GTECH_XNOR2 U430 ( .A(n340), .B(n11), .Z(n458) );
  GTECH_NOT U431 ( .A(n459), .Z(n457) );
  GTECH_OAI21 U432 ( .A(n12), .B(n455), .C(n460), .Z(N135) );
  GTECH_OAI21 U433 ( .A(n388), .B(n384), .C(n366), .Z(n460) );
  GTECH_OAI21 U434 ( .A(n12), .B(n461), .C(n454), .Z(n366) );
  GTECH_NOT U435 ( .A(n462), .Z(n384) );
  GTECH_NAND3 U436 ( .A(n28), .B(n463), .C(N155), .Z(n462) );
  GTECH_NOT U437 ( .A(n464), .Z(n388) );
  GTECH_NAND3 U438 ( .A(n10), .B(n465), .C(N155), .Z(n464) );
  GTECH_NAND2 U439 ( .A(n466), .B(N155), .Z(n455) );
  GTECH_XNOR2 U440 ( .A(n28), .B(n10), .Z(n466) );
  GTECH_AND2 U441 ( .A(N155), .B(n467), .Z(N134) );
  GTECH_NOT U442 ( .A(n13), .Z(n467) );
  GTECH_AND2 U443 ( .A(N155), .B(n468), .Z(N133) );
  GTECH_NOT U444 ( .A(n14), .Z(n468) );
  GTECH_AND2 U445 ( .A(N155), .B(n469), .Z(N132) );
  GTECH_NOT U446 ( .A(n15), .Z(n469) );
  GTECH_AND2 U447 ( .A(N155), .B(n470), .Z(N131) );
  GTECH_NOT U448 ( .A(n16), .Z(n470) );
  GTECH_AND2 U449 ( .A(N155), .B(n471), .Z(N130) );
  GTECH_NOT U450 ( .A(n17), .Z(n471) );
  GTECH_AND2 U451 ( .A(N155), .B(n472), .Z(N129) );
  GTECH_NOT U452 ( .A(n18), .Z(n472) );
  GTECH_AND2 U453 ( .A(N155), .B(n473), .Z(N128) );
  GTECH_NOT U454 ( .A(n19), .Z(n473) );
  GTECH_AND2 U455 ( .A(N155), .B(n474), .Z(N127) );
  GTECH_NOT U456 ( .A(n20), .Z(n474) );
  GTECH_AND2 U457 ( .A(N155), .B(n475), .Z(N126) );
  GTECH_NOT U458 ( .A(n21), .Z(n475) );
  GTECH_AND2 U459 ( .A(N155), .B(n476), .Z(N125) );
  GTECH_NOT U460 ( .A(n22), .Z(n476) );
  GTECH_AND2 U461 ( .A(N155), .B(n477), .Z(N124) );
  GTECH_NOT U462 ( .A(n23), .Z(n477) );
  GTECH_AND2 U463 ( .A(N155), .B(n478), .Z(N123) );
  GTECH_NOT U464 ( .A(n24), .Z(n478) );
  GTECH_AND2 U465 ( .A(N155), .B(n479), .Z(N122) );
  GTECH_NOT U466 ( .A(n25), .Z(n479) );
  GTECH_AND2 U467 ( .A(N155), .B(n480), .Z(N121) );
  GTECH_NOT U468 ( .A(n26), .Z(n480) );
  GTECH_AND2 U469 ( .A(N155), .B(n481), .Z(N120) );
  GTECH_NOT U470 ( .A(n27), .Z(n481) );
  GTECH_NOT U471 ( .A(n390), .Z(N155) );
  GTECH_NAND4 U472 ( .A(n8), .B(n7), .C(n9), .D(n482), .Z(n390) );
  GTECH_AND3 U473 ( .A(n377), .B(n396), .C(n6), .Z(n482) );
  GTECH_NOT U474 ( .A(n338), .Z(n396) );
  GTECH_NOT U475 ( .A(n483), .Z(N116) );
  GTECH_AOI222 U476 ( .A(n359), .B(n387), .C(n361), .D(n389), .E(n385), .F(
        n357), .Z(n483) );
  GTECH_XNOR2 U477 ( .A(n484), .B(n485), .Z(n385) );
  GTECH_NOT U478 ( .A(n486), .Z(n485) );
  GTECH_ADD_ABC U479 ( .A(n354), .B(n31), .C(n487), .COUT(n484) );
  GTECH_XNOR2 U480 ( .A(n488), .B(n486), .Z(n389) );
  GTECH_XNOR2 U481 ( .A(n355), .B(n30), .Z(n486) );
  GTECH_AND2 U482 ( .A(n489), .B(n490), .Z(n488) );
  GTECH_OAI21 U483 ( .A(n354), .B(n393), .C(n491), .Z(n490) );
  GTECH_OR_NOT U484 ( .A(n31), .B(n354), .Z(n489) );
  GTECH_NOT U485 ( .A(n30), .Z(n387) );
  GTECH_NAND2 U486 ( .A(n370), .B(n492), .Z(N115) );
  GTECH_NOT U487 ( .A(N41), .Z(n492) );
  GTECH_NAND2 U488 ( .A(n377), .B(n371), .Z(N41) );
  GTECH_NAND2 U489 ( .A(Ld), .B(n377), .Z(n371) );
  GTECH_NOT U490 ( .A(n493), .Z(N113) );
  GTECH_AOI222 U491 ( .A(n359), .B(n393), .C(n361), .D(n394), .E(n392), .F(
        n357), .Z(n493) );
  GTECH_XNOR2 U492 ( .A(n487), .B(n494), .Z(n392) );
  GTECH_ADD_ABC U493 ( .A(n353), .B(n32), .C(n495), .COUT(n487) );
  GTECH_NOT U494 ( .A(n496), .Z(n394) );
  GTECH_XNOR2 U495 ( .A(n497), .B(n494), .Z(n496) );
  GTECH_NOT U496 ( .A(n498), .Z(n494) );
  GTECH_XNOR2 U497 ( .A(n354), .B(n31), .Z(n498) );
  GTECH_NOT U498 ( .A(n491), .Z(n497) );
  GTECH_OAI21 U499 ( .A(n32), .B(n499), .C(n500), .Z(n491) );
  GTECH_OAI21 U500 ( .A(n353), .B(n399), .C(n501), .Z(n500) );
  GTECH_NOT U501 ( .A(n353), .Z(n499) );
  GTECH_NOT U502 ( .A(n31), .Z(n393) );
  GTECH_NOT U503 ( .A(n502), .Z(N112) );
  GTECH_AOI222 U504 ( .A(n359), .B(n399), .C(n361), .D(n400), .E(n398), .F(
        n357), .Z(n502) );
  GTECH_XNOR2 U505 ( .A(n495), .B(n503), .Z(n398) );
  GTECH_ADD_ABC U506 ( .A(n33), .B(n352), .C(n504), .COUT(n495) );
  GTECH_NOT U507 ( .A(n505), .Z(n400) );
  GTECH_XNOR2 U508 ( .A(n506), .B(n503), .Z(n505) );
  GTECH_NOT U509 ( .A(n507), .Z(n503) );
  GTECH_XNOR2 U510 ( .A(n353), .B(n32), .Z(n507) );
  GTECH_NOT U511 ( .A(n501), .Z(n506) );
  GTECH_OAI21 U512 ( .A(n33), .B(n508), .C(n509), .Z(n501) );
  GTECH_OAI21 U513 ( .A(n352), .B(n403), .C(n510), .Z(n509) );
  GTECH_NOT U514 ( .A(n352), .Z(n508) );
  GTECH_NOT U515 ( .A(n32), .Z(n399) );
  GTECH_NOT U516 ( .A(n511), .Z(N111) );
  GTECH_AOI222 U517 ( .A(n359), .B(n403), .C(n361), .D(n404), .E(n402), .F(
        n357), .Z(n511) );
  GTECH_XNOR2 U518 ( .A(n504), .B(n512), .Z(n402) );
  GTECH_ADD_ABC U519 ( .A(n34), .B(n351), .C(n513), .COUT(n504) );
  GTECH_NOT U520 ( .A(n514), .Z(n404) );
  GTECH_XNOR2 U521 ( .A(n515), .B(n512), .Z(n514) );
  GTECH_NOT U522 ( .A(n516), .Z(n512) );
  GTECH_XNOR2 U523 ( .A(n33), .B(n352), .Z(n516) );
  GTECH_NOT U524 ( .A(n510), .Z(n515) );
  GTECH_OAI21 U525 ( .A(n34), .B(n517), .C(n518), .Z(n510) );
  GTECH_OAI21 U526 ( .A(n351), .B(n407), .C(n519), .Z(n518) );
  GTECH_NOT U527 ( .A(n351), .Z(n517) );
  GTECH_NOT U528 ( .A(n33), .Z(n403) );
  GTECH_NOT U529 ( .A(n520), .Z(N110) );
  GTECH_AOI222 U530 ( .A(n359), .B(n407), .C(n361), .D(n408), .E(n406), .F(
        n357), .Z(n520) );
  GTECH_XNOR2 U531 ( .A(n513), .B(n521), .Z(n406) );
  GTECH_ADD_ABC U532 ( .A(n35), .B(n350), .C(n522), .COUT(n513) );
  GTECH_NOT U533 ( .A(n523), .Z(n408) );
  GTECH_XNOR2 U534 ( .A(n524), .B(n521), .Z(n523) );
  GTECH_NOT U535 ( .A(n525), .Z(n521) );
  GTECH_XNOR2 U536 ( .A(n34), .B(n351), .Z(n525) );
  GTECH_NOT U537 ( .A(n519), .Z(n524) );
  GTECH_OAI21 U538 ( .A(n35), .B(n526), .C(n527), .Z(n519) );
  GTECH_OAI21 U539 ( .A(n350), .B(n411), .C(n528), .Z(n527) );
  GTECH_NOT U540 ( .A(n350), .Z(n526) );
  GTECH_NOT U541 ( .A(n34), .Z(n407) );
  GTECH_NOT U542 ( .A(n529), .Z(N109) );
  GTECH_AOI222 U543 ( .A(n359), .B(n411), .C(n361), .D(n412), .E(n410), .F(
        n357), .Z(n529) );
  GTECH_XNOR2 U544 ( .A(n522), .B(n530), .Z(n410) );
  GTECH_ADD_ABC U545 ( .A(n36), .B(n349), .C(n531), .COUT(n522) );
  GTECH_NOT U546 ( .A(n532), .Z(n412) );
  GTECH_XNOR2 U547 ( .A(n533), .B(n530), .Z(n532) );
  GTECH_NOT U548 ( .A(n534), .Z(n530) );
  GTECH_XNOR2 U549 ( .A(n35), .B(n350), .Z(n534) );
  GTECH_NOT U550 ( .A(n528), .Z(n533) );
  GTECH_OAI21 U551 ( .A(n36), .B(n535), .C(n536), .Z(n528) );
  GTECH_OAI21 U552 ( .A(n349), .B(n415), .C(n537), .Z(n536) );
  GTECH_NOT U553 ( .A(n349), .Z(n535) );
  GTECH_NOT U554 ( .A(n35), .Z(n411) );
  GTECH_NOT U555 ( .A(n538), .Z(N108) );
  GTECH_AOI222 U556 ( .A(n359), .B(n415), .C(n361), .D(n416), .E(n414), .F(
        n357), .Z(n538) );
  GTECH_XNOR2 U557 ( .A(n531), .B(n539), .Z(n414) );
  GTECH_ADD_ABC U558 ( .A(n37), .B(n348), .C(n540), .COUT(n531) );
  GTECH_NOT U559 ( .A(n541), .Z(n416) );
  GTECH_XNOR2 U560 ( .A(n542), .B(n539), .Z(n541) );
  GTECH_NOT U561 ( .A(n543), .Z(n539) );
  GTECH_XNOR2 U562 ( .A(n36), .B(n349), .Z(n543) );
  GTECH_NOT U563 ( .A(n537), .Z(n542) );
  GTECH_OAI21 U564 ( .A(n37), .B(n544), .C(n545), .Z(n537) );
  GTECH_OAI21 U565 ( .A(n348), .B(n419), .C(n546), .Z(n545) );
  GTECH_NOT U566 ( .A(n348), .Z(n544) );
  GTECH_NOT U567 ( .A(n36), .Z(n415) );
  GTECH_NOT U568 ( .A(n547), .Z(N107) );
  GTECH_AOI222 U569 ( .A(n359), .B(n419), .C(n361), .D(n420), .E(n418), .F(
        n357), .Z(n547) );
  GTECH_XNOR2 U570 ( .A(n540), .B(n548), .Z(n418) );
  GTECH_ADD_ABC U571 ( .A(n38), .B(n347), .C(n549), .COUT(n540) );
  GTECH_NOT U572 ( .A(n550), .Z(n420) );
  GTECH_XNOR2 U573 ( .A(n551), .B(n548), .Z(n550) );
  GTECH_NOT U574 ( .A(n552), .Z(n548) );
  GTECH_XNOR2 U575 ( .A(n37), .B(n348), .Z(n552) );
  GTECH_NOT U576 ( .A(n546), .Z(n551) );
  GTECH_OAI21 U577 ( .A(n38), .B(n553), .C(n554), .Z(n546) );
  GTECH_OAI21 U578 ( .A(n347), .B(n423), .C(n555), .Z(n554) );
  GTECH_NOT U579 ( .A(n347), .Z(n553) );
  GTECH_NOT U580 ( .A(n37), .Z(n419) );
  GTECH_NOT U581 ( .A(n556), .Z(N106) );
  GTECH_AOI222 U582 ( .A(n359), .B(n423), .C(n361), .D(n424), .E(n422), .F(
        n357), .Z(n556) );
  GTECH_XNOR2 U583 ( .A(n549), .B(n557), .Z(n422) );
  GTECH_ADD_ABC U584 ( .A(n39), .B(n346), .C(n558), .COUT(n549) );
  GTECH_NOT U585 ( .A(n559), .Z(n424) );
  GTECH_XNOR2 U586 ( .A(n560), .B(n557), .Z(n559) );
  GTECH_NOT U587 ( .A(n561), .Z(n557) );
  GTECH_XNOR2 U588 ( .A(n38), .B(n347), .Z(n561) );
  GTECH_NOT U589 ( .A(n555), .Z(n560) );
  GTECH_OAI21 U590 ( .A(n39), .B(n562), .C(n563), .Z(n555) );
  GTECH_OAI21 U591 ( .A(n346), .B(n427), .C(n564), .Z(n563) );
  GTECH_NOT U592 ( .A(n346), .Z(n562) );
  GTECH_NOT U593 ( .A(n38), .Z(n423) );
  GTECH_NOT U594 ( .A(n565), .Z(N105) );
  GTECH_AOI222 U595 ( .A(n359), .B(n427), .C(n361), .D(n428), .E(n426), .F(
        n357), .Z(n565) );
  GTECH_XNOR2 U596 ( .A(n558), .B(n566), .Z(n426) );
  GTECH_ADD_ABC U597 ( .A(n40), .B(n345), .C(n567), .COUT(n558) );
  GTECH_NOT U598 ( .A(n568), .Z(n428) );
  GTECH_XNOR2 U599 ( .A(n569), .B(n566), .Z(n568) );
  GTECH_NOT U600 ( .A(n570), .Z(n566) );
  GTECH_XNOR2 U601 ( .A(n39), .B(n346), .Z(n570) );
  GTECH_NOT U602 ( .A(n564), .Z(n569) );
  GTECH_OAI21 U603 ( .A(n40), .B(n571), .C(n572), .Z(n564) );
  GTECH_OAI21 U604 ( .A(n345), .B(n431), .C(n573), .Z(n572) );
  GTECH_NOT U605 ( .A(n345), .Z(n571) );
  GTECH_NOT U606 ( .A(n39), .Z(n427) );
  GTECH_NOT U607 ( .A(n574), .Z(N104) );
  GTECH_AOI222 U608 ( .A(n359), .B(n431), .C(n361), .D(n432), .E(n430), .F(
        n357), .Z(n574) );
  GTECH_XNOR2 U609 ( .A(n567), .B(n575), .Z(n430) );
  GTECH_ADD_ABC U610 ( .A(n41), .B(n344), .C(n576), .COUT(n567) );
  GTECH_NOT U611 ( .A(n577), .Z(n432) );
  GTECH_XNOR2 U612 ( .A(n578), .B(n575), .Z(n577) );
  GTECH_NOT U613 ( .A(n579), .Z(n575) );
  GTECH_XNOR2 U614 ( .A(n40), .B(n345), .Z(n579) );
  GTECH_NOT U615 ( .A(n573), .Z(n578) );
  GTECH_OAI21 U616 ( .A(n41), .B(n580), .C(n581), .Z(n573) );
  GTECH_OAI21 U617 ( .A(n344), .B(n435), .C(n582), .Z(n581) );
  GTECH_NOT U618 ( .A(n344), .Z(n580) );
  GTECH_NOT U619 ( .A(n40), .Z(n431) );
  GTECH_NOT U620 ( .A(n583), .Z(N103) );
  GTECH_AOI222 U621 ( .A(n359), .B(n435), .C(n361), .D(n436), .E(n434), .F(
        n357), .Z(n583) );
  GTECH_XNOR2 U622 ( .A(n576), .B(n584), .Z(n434) );
  GTECH_ADD_ABC U623 ( .A(n42), .B(n343), .C(n585), .COUT(n576) );
  GTECH_NOT U624 ( .A(n586), .Z(n436) );
  GTECH_XNOR2 U625 ( .A(n587), .B(n584), .Z(n586) );
  GTECH_NOT U626 ( .A(n588), .Z(n584) );
  GTECH_XNOR2 U627 ( .A(n41), .B(n344), .Z(n588) );
  GTECH_NOT U628 ( .A(n582), .Z(n587) );
  GTECH_OAI21 U629 ( .A(n42), .B(n589), .C(n590), .Z(n582) );
  GTECH_OAI21 U630 ( .A(n343), .B(n440), .C(n591), .Z(n590) );
  GTECH_NOT U631 ( .A(n343), .Z(n589) );
  GTECH_NOT U632 ( .A(n41), .Z(n435) );
  GTECH_NOT U633 ( .A(n592), .Z(N102) );
  GTECH_AOI222 U634 ( .A(n359), .B(n440), .C(n361), .D(n441), .E(n439), .F(
        n357), .Z(n592) );
  GTECH_XNOR2 U635 ( .A(n585), .B(n593), .Z(n439) );
  GTECH_ADD_ABC U636 ( .A(n43), .B(n342), .C(n594), .COUT(n585) );
  GTECH_NOT U637 ( .A(n595), .Z(n441) );
  GTECH_XNOR2 U638 ( .A(n596), .B(n593), .Z(n595) );
  GTECH_NOT U639 ( .A(n597), .Z(n593) );
  GTECH_XNOR2 U640 ( .A(n42), .B(n343), .Z(n597) );
  GTECH_NOT U641 ( .A(n591), .Z(n596) );
  GTECH_OAI21 U642 ( .A(n43), .B(n598), .C(n599), .Z(n591) );
  GTECH_OAI21 U643 ( .A(n342), .B(n444), .C(n600), .Z(n599) );
  GTECH_NOT U644 ( .A(n342), .Z(n598) );
  GTECH_NOT U645 ( .A(n42), .Z(n440) );
  GTECH_NOT U646 ( .A(n601), .Z(N101) );
  GTECH_AOI222 U647 ( .A(n359), .B(n444), .C(n361), .D(n445), .E(n443), .F(
        n357), .Z(n601) );
  GTECH_XNOR2 U648 ( .A(n594), .B(n602), .Z(n443) );
  GTECH_ADD_ABC U649 ( .A(n29), .B(n341), .C(n603), .COUT(n594) );
  GTECH_NOT U650 ( .A(n604), .Z(n445) );
  GTECH_XNOR2 U651 ( .A(n605), .B(n602), .Z(n604) );
  GTECH_NOT U652 ( .A(n606), .Z(n602) );
  GTECH_XNOR2 U653 ( .A(n43), .B(n342), .Z(n606) );
  GTECH_NOT U654 ( .A(n600), .Z(n605) );
  GTECH_OAI21 U655 ( .A(n29), .B(n607), .C(n608), .Z(n600) );
  GTECH_OAI21 U656 ( .A(n341), .B(n448), .C(n609), .Z(n608) );
  GTECH_NOT U657 ( .A(n341), .Z(n607) );
  GTECH_NOT U658 ( .A(n43), .Z(n444) );
  GTECH_NOT U659 ( .A(n610), .Z(N100) );
  GTECH_AOI222 U660 ( .A(n447), .B(n357), .C(n359), .D(n448), .E(n361), .F(
        n449), .Z(n610) );
  GTECH_NOT U661 ( .A(n611), .Z(n449) );
  GTECH_XNOR2 U662 ( .A(n612), .B(n613), .Z(n611) );
  GTECH_NOT U663 ( .A(n609), .Z(n612) );
  GTECH_OAI21 U664 ( .A(n11), .B(n614), .C(n615), .Z(n609) );
  GTECH_OAI21 U665 ( .A(n340), .B(n360), .C(n454), .Z(n615) );
  GTECH_NAND2 U666 ( .A(n12), .B(n461), .Z(n454) );
  GTECH_NOT U667 ( .A(n11), .Z(n360) );
  GTECH_NOT U668 ( .A(n340), .Z(n614) );
  GTECH_NOT U669 ( .A(n369), .Z(n361) );
  GTECH_NAND2 U670 ( .A(N82), .B(n10), .Z(n369) );
  GTECH_NOT U671 ( .A(n616), .Z(N82) );
  GTECH_NOT U672 ( .A(n29), .Z(n448) );
  GTECH_NOT U673 ( .A(n617), .Z(n359) );
  GTECH_MUX2 U674 ( .A(n616), .B(n618), .S(n10), .Z(n617) );
  GTECH_NAND2 U675 ( .A(n28), .B(n375), .Z(n618) );
  GTECH_NAND2 U676 ( .A(n375), .B(n465), .Z(n616) );
  GTECH_NOT U677 ( .A(n28), .Z(n465) );
  GTECH_NOT U678 ( .A(n368), .Z(n357) );
  GTECH_NAND3 U679 ( .A(n375), .B(n463), .C(n28), .Z(n368) );
  GTECH_NOT U680 ( .A(n10), .Z(n463) );
  GTECH_NOT U681 ( .A(n370), .Z(n375) );
  GTECH_OAI21 U682 ( .A(n373), .B(n374), .C(n619), .Z(n370) );
  GTECH_AND2 U683 ( .A(n376), .B(n377), .Z(n619) );
  GTECH_NOT U684 ( .A(Rst), .Z(n377) );
  GTECH_NOT U685 ( .A(Ld), .Z(n376) );
  GTECH_NOT U686 ( .A(n9), .Z(n374) );
  GTECH_NAND2 U687 ( .A(n8), .B(n379), .Z(n373) );
  GTECH_NOT U688 ( .A(n382), .Z(n379) );
  GTECH_NAND2 U689 ( .A(n7), .B(n381), .Z(n382) );
  GTECH_NOT U690 ( .A(n620), .Z(n381) );
  GTECH_NAND2 U691 ( .A(n6), .B(n338), .Z(n620) );
  GTECH_XNOR2 U692 ( .A(n603), .B(n613), .Z(n447) );
  GTECH_NOT U693 ( .A(n621), .Z(n613) );
  GTECH_XNOR2 U694 ( .A(n29), .B(n341), .Z(n621) );
  GTECH_ADD_ABC U695 ( .A(n340), .B(n11), .C(n459), .COUT(n603) );
  GTECH_NAND2 U696 ( .A(n364), .B(n461), .Z(n459) );
  GTECH_NOT U697 ( .A(n339), .Z(n461) );
  GTECH_NOT U698 ( .A(n12), .Z(n364) );
endmodule

