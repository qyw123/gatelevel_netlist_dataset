
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392;

  GTECH_MUX2 U142 ( .A(n281), .B(n282), .S(n283), .Z(sum[9]) );
  GTECH_XOR2 U143 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_XOR2 U144 ( .A(n286), .B(n285), .Z(n281) );
  GTECH_AOI21 U145 ( .A(n287), .B(n288), .C(n289), .Z(n285) );
  GTECH_NOT U146 ( .A(b[9]), .Z(n288) );
  GTECH_XOR2 U147 ( .A(n290), .B(n283), .Z(sum[8]) );
  GTECH_MUX2 U148 ( .A(n291), .B(n292), .S(n293), .Z(sum[7]) );
  GTECH_XOR2 U149 ( .A(n294), .B(n295), .Z(n292) );
  GTECH_XNOR2 U150 ( .A(n294), .B(n296), .Z(n291) );
  GTECH_AND2 U151 ( .A(n297), .B(n298), .Z(n296) );
  GTECH_OAI21 U152 ( .A(b[6]), .B(a[6]), .C(n299), .Z(n298) );
  GTECH_XOR2 U153 ( .A(a[7]), .B(b[7]), .Z(n294) );
  GTECH_OAI21 U154 ( .A(n300), .B(n297), .C(n301), .Z(sum[6]) );
  GTECH_MUX2 U155 ( .A(n302), .B(n303), .S(b[6]), .Z(n301) );
  GTECH_OR_NOT U156 ( .A(a[6]), .B(n300), .Z(n303) );
  GTECH_XNOR2 U157 ( .A(n304), .B(n300), .Z(n302) );
  GTECH_NOT U158 ( .A(a[6]), .Z(n304) );
  GTECH_AOI21 U159 ( .A(n305), .B(n293), .C(n299), .Z(n300) );
  GTECH_OAI21 U160 ( .A(n306), .B(n307), .C(n308), .Z(n299) );
  GTECH_MUX2 U161 ( .A(n309), .B(n310), .S(n311), .Z(sum[5]) );
  GTECH_AND2 U162 ( .A(n308), .B(n312), .Z(n311) );
  GTECH_OAI21 U163 ( .A(a[4]), .B(n293), .C(n313), .Z(n310) );
  GTECH_OAI21 U164 ( .A(n314), .B(n315), .C(n316), .Z(n313) );
  GTECH_OAI21 U165 ( .A(n317), .B(n314), .C(n307), .Z(n309) );
  GTECH_OR_NOT U166 ( .A(n316), .B(a[4]), .Z(n307) );
  GTECH_XOR2 U167 ( .A(n318), .B(n314), .Z(sum[4]) );
  GTECH_NOT U168 ( .A(n293), .Z(n314) );
  GTECH_MUX2 U169 ( .A(n319), .B(n320), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U170 ( .A(n321), .B(n322), .Z(n320) );
  GTECH_XOR2 U171 ( .A(n323), .B(n321), .Z(n319) );
  GTECH_XOR2 U172 ( .A(a[3]), .B(b[3]), .Z(n321) );
  GTECH_AOI21 U173 ( .A(n324), .B(n325), .C(n326), .Z(n323) );
  GTECH_OA21 U174 ( .A(n325), .B(n324), .C(n327), .Z(n326) );
  GTECH_MUX2 U175 ( .A(n328), .B(n329), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U176 ( .A(n330), .B(n331), .Z(n329) );
  GTECH_XOR2 U177 ( .A(n330), .B(n325), .Z(n328) );
  GTECH_AOI21 U178 ( .A(n332), .B(n333), .C(n334), .Z(n325) );
  GTECH_XNOR2 U179 ( .A(n324), .B(n327), .Z(n330) );
  GTECH_NOT U180 ( .A(b[2]), .Z(n327) );
  GTECH_MUX2 U181 ( .A(n335), .B(n336), .S(n337), .Z(sum[1]) );
  GTECH_AND_NOT U182 ( .A(n332), .B(n334), .Z(n337) );
  GTECH_OAI21 U183 ( .A(cin), .B(n333), .C(n338), .Z(n336) );
  GTECH_NOT U184 ( .A(n339), .Z(n335) );
  GTECH_AOI21 U185 ( .A(n338), .B(cin), .C(n333), .Z(n339) );
  GTECH_MUX2 U186 ( .A(n340), .B(n341), .S(n342), .Z(sum[15]) );
  GTECH_XOR2 U187 ( .A(n343), .B(n344), .Z(n341) );
  GTECH_AND2 U188 ( .A(n345), .B(n346), .Z(n344) );
  GTECH_OAI21 U189 ( .A(b[14]), .B(a[14]), .C(n347), .Z(n345) );
  GTECH_XNOR2 U190 ( .A(n343), .B(n348), .Z(n340) );
  GTECH_XNOR2 U191 ( .A(a[15]), .B(b[15]), .Z(n343) );
  GTECH_OAI21 U192 ( .A(n349), .B(n346), .C(n350), .Z(sum[14]) );
  GTECH_MUX2 U193 ( .A(n351), .B(n352), .S(b[14]), .Z(n350) );
  GTECH_OR_NOT U194 ( .A(a[14]), .B(n349), .Z(n352) );
  GTECH_XNOR2 U195 ( .A(n353), .B(n349), .Z(n351) );
  GTECH_AOI21 U196 ( .A(n354), .B(n355), .C(n347), .Z(n349) );
  GTECH_OAI2N2 U197 ( .A(n356), .B(n357), .C(a[13]), .D(b[13]), .Z(n347) );
  GTECH_NOT U198 ( .A(n342), .Z(n355) );
  GTECH_MUX2 U199 ( .A(n358), .B(n359), .S(n342), .Z(sum[13]) );
  GTECH_XNOR2 U200 ( .A(n357), .B(n360), .Z(n359) );
  GTECH_XOR2 U201 ( .A(n361), .B(n360), .Z(n358) );
  GTECH_AOI21 U202 ( .A(a[13]), .B(b[13]), .C(n356), .Z(n360) );
  GTECH_NOT U203 ( .A(n362), .Z(n356) );
  GTECH_OR_NOT U204 ( .A(n363), .B(n364), .Z(sum[12]) );
  GTECH_AOI21 U205 ( .A(n357), .B(n361), .C(n342), .Z(n363) );
  GTECH_MUX2 U206 ( .A(n365), .B(n366), .S(n283), .Z(sum[11]) );
  GTECH_XNOR2 U207 ( .A(n367), .B(n368), .Z(n366) );
  GTECH_OA21 U208 ( .A(n369), .B(n370), .C(n371), .Z(n368) );
  GTECH_XOR2 U209 ( .A(n367), .B(n372), .Z(n365) );
  GTECH_XOR2 U210 ( .A(a[11]), .B(b[11]), .Z(n367) );
  GTECH_MUX2 U211 ( .A(n373), .B(n374), .S(n375), .Z(sum[10]) );
  GTECH_OA21 U212 ( .A(n283), .B(n376), .C(n370), .Z(n375) );
  GTECH_OAI21 U213 ( .A(n284), .B(n289), .C(n377), .Z(n370) );
  GTECH_XOR2 U214 ( .A(b[10]), .B(a[10]), .Z(n374) );
  GTECH_OR_NOT U215 ( .A(n369), .B(n371), .Z(n373) );
  GTECH_XOR2 U216 ( .A(cin), .B(n378), .Z(sum[0]) );
  GTECH_OAI21 U217 ( .A(n379), .B(n342), .C(n364), .Z(cout) );
  GTECH_NAND3 U218 ( .A(n361), .B(n357), .C(n342), .Z(n364) );
  GTECH_NAND2 U219 ( .A(b[12]), .B(a[12]), .Z(n357) );
  GTECH_MUX2 U220 ( .A(n380), .B(n290), .S(n283), .Z(n342) );
  GTECH_MUX2 U221 ( .A(n318), .B(n381), .S(n293), .Z(n283) );
  GTECH_MUX2 U222 ( .A(n378), .B(n382), .S(cin), .Z(n293) );
  GTECH_OA21 U223 ( .A(a[3]), .B(n322), .C(n383), .Z(n382) );
  GTECH_NOT U224 ( .A(n384), .Z(n383) );
  GTECH_AOI21 U225 ( .A(n322), .B(a[3]), .C(b[3]), .Z(n384) );
  GTECH_OAI21 U226 ( .A(n385), .B(n324), .C(n386), .Z(n322) );
  GTECH_OAI21 U227 ( .A(a[2]), .B(n331), .C(b[2]), .Z(n386) );
  GTECH_NOT U228 ( .A(n385), .Z(n331) );
  GTECH_NOT U229 ( .A(a[2]), .Z(n324) );
  GTECH_AOI21 U230 ( .A(n332), .B(n338), .C(n334), .Z(n385) );
  GTECH_AND2 U231 ( .A(b[1]), .B(a[1]), .Z(n334) );
  GTECH_OR2 U232 ( .A(a[1]), .B(b[1]), .Z(n332) );
  GTECH_AND_NOT U233 ( .A(n338), .B(n333), .Z(n378) );
  GTECH_AND2 U234 ( .A(b[0]), .B(a[0]), .Z(n333) );
  GTECH_OR2 U235 ( .A(b[0]), .B(a[0]), .Z(n338) );
  GTECH_AOI21 U236 ( .A(n295), .B(a[7]), .C(n387), .Z(n381) );
  GTECH_OA21 U237 ( .A(a[7]), .B(n295), .C(b[7]), .Z(n387) );
  GTECH_NAND2 U238 ( .A(n388), .B(n297), .Z(n295) );
  GTECH_NAND2 U239 ( .A(a[6]), .B(b[6]), .Z(n297) );
  GTECH_OAI21 U240 ( .A(a[6]), .B(b[6]), .C(n305), .Z(n388) );
  GTECH_OAI21 U241 ( .A(n317), .B(n306), .C(n308), .Z(n305) );
  GTECH_NAND2 U242 ( .A(a[5]), .B(b[5]), .Z(n308) );
  GTECH_NOT U243 ( .A(n312), .Z(n306) );
  GTECH_OR2 U244 ( .A(a[5]), .B(b[5]), .Z(n312) );
  GTECH_AND2 U245 ( .A(n315), .B(n316), .Z(n317) );
  GTECH_NOT U246 ( .A(a[4]), .Z(n315) );
  GTECH_XOR2 U247 ( .A(a[4]), .B(n316), .Z(n318) );
  GTECH_NOT U248 ( .A(b[4]), .Z(n316) );
  GTECH_OR_NOT U249 ( .A(n284), .B(n286), .Z(n290) );
  GTECH_AND2 U250 ( .A(b[8]), .B(a[8]), .Z(n284) );
  GTECH_AOI21 U251 ( .A(n372), .B(a[11]), .C(n389), .Z(n380) );
  GTECH_OA21 U252 ( .A(a[11]), .B(n372), .C(b[11]), .Z(n389) );
  GTECH_OAI21 U253 ( .A(n369), .B(n376), .C(n371), .Z(n372) );
  GTECH_NAND2 U254 ( .A(a[10]), .B(b[10]), .Z(n371) );
  GTECH_OAI21 U255 ( .A(n289), .B(n286), .C(n377), .Z(n376) );
  GTECH_OR_NOT U256 ( .A(b[9]), .B(n287), .Z(n377) );
  GTECH_NOT U257 ( .A(a[9]), .Z(n287) );
  GTECH_OR2 U258 ( .A(a[8]), .B(b[8]), .Z(n286) );
  GTECH_AND2 U259 ( .A(a[9]), .B(b[9]), .Z(n289) );
  GTECH_AND_NOT U260 ( .A(n390), .B(b[10]), .Z(n369) );
  GTECH_NOT U261 ( .A(a[10]), .Z(n390) );
  GTECH_AOI21 U262 ( .A(n348), .B(a[15]), .C(n391), .Z(n379) );
  GTECH_OA21 U263 ( .A(a[15]), .B(n348), .C(b[15]), .Z(n391) );
  GTECH_NAND2 U264 ( .A(n392), .B(n346), .Z(n348) );
  GTECH_OR_NOT U265 ( .A(n353), .B(b[14]), .Z(n346) );
  GTECH_NOT U266 ( .A(a[14]), .Z(n353) );
  GTECH_OAI21 U267 ( .A(a[14]), .B(b[14]), .C(n354), .Z(n392) );
  GTECH_AO22 U268 ( .A(a[13]), .B(b[13]), .C(n362), .D(n361), .Z(n354) );
  GTECH_OR2 U269 ( .A(a[12]), .B(b[12]), .Z(n361) );
  GTECH_OR2 U270 ( .A(b[13]), .B(a[13]), .Z(n362) );
endmodule

