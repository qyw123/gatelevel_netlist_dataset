
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377;

  GTECH_OAI22 U131 ( .A(n270), .B(n271), .C(n272), .D(n273), .Z(sum[9]) );
  GTECH_XOR2 U132 ( .A(n274), .B(n275), .Z(n273) );
  GTECH_XNOR2 U133 ( .A(n275), .B(n276), .Z(n270) );
  GTECH_NOT U134 ( .A(n277), .Z(n276) );
  GTECH_OAI21 U135 ( .A(a[9]), .B(b[9]), .C(n278), .Z(n275) );
  GTECH_OAI21 U136 ( .A(n279), .B(n271), .C(n280), .Z(sum[8]) );
  GTECH_OAI22 U137 ( .A(n281), .B(n282), .C(n283), .D(n284), .Z(sum[7]) );
  GTECH_XNOR2 U138 ( .A(n285), .B(n286), .Z(n283) );
  GTECH_XNOR2 U139 ( .A(n286), .B(n287), .Z(n282) );
  GTECH_AOI21 U140 ( .A(n288), .B(n289), .C(n290), .Z(n287) );
  GTECH_AOI21 U141 ( .A(n291), .B(a[6]), .C(b[6]), .Z(n290) );
  GTECH_XOR2 U142 ( .A(a[7]), .B(b[7]), .Z(n286) );
  GTECH_OAI22 U143 ( .A(n292), .B(n281), .C(n293), .D(n284), .Z(sum[6]) );
  GTECH_XOR2 U144 ( .A(n294), .B(n295), .Z(n293) );
  GTECH_XNOR2 U145 ( .A(n291), .B(n295), .Z(n292) );
  GTECH_XOR2 U146 ( .A(a[6]), .B(b[6]), .Z(n295) );
  GTECH_NOT U147 ( .A(n289), .Z(n291) );
  GTECH_OA21 U148 ( .A(n296), .B(n297), .C(n298), .Z(n289) );
  GTECH_OAI2N2 U149 ( .A(n299), .B(n300), .C(n300), .D(n301), .Z(sum[5]) );
  GTECH_NOT U150 ( .A(n302), .Z(n301) );
  GTECH_OA21 U151 ( .A(n303), .B(n284), .C(n297), .Z(n302) );
  GTECH_OR_NOT U152 ( .A(n304), .B(b[4]), .Z(n297) );
  GTECH_OR_NOT U153 ( .A(n296), .B(n298), .Z(n300) );
  GTECH_AOI21 U154 ( .A(n304), .B(n284), .C(n305), .Z(n299) );
  GTECH_AOI21 U155 ( .A(n281), .B(a[4]), .C(b[4]), .Z(n305) );
  GTECH_NOT U156 ( .A(n284), .Z(n281) );
  GTECH_XOR2 U157 ( .A(n306), .B(n284), .Z(sum[4]) );
  GTECH_OAI22 U158 ( .A(n307), .B(n308), .C(cin), .D(n309), .Z(sum[3]) );
  GTECH_XNOR2 U159 ( .A(n310), .B(n311), .Z(n309) );
  GTECH_AOI21 U160 ( .A(n312), .B(n313), .C(n314), .Z(n311) );
  GTECH_AOI21 U161 ( .A(n315), .B(a[2]), .C(b[2]), .Z(n314) );
  GTECH_NOT U162 ( .A(n313), .Z(n315) );
  GTECH_XNOR2 U163 ( .A(n316), .B(n310), .Z(n308) );
  GTECH_XOR2 U164 ( .A(a[3]), .B(b[3]), .Z(n310) );
  GTECH_OAI22 U165 ( .A(n307), .B(n317), .C(cin), .D(n318), .Z(sum[2]) );
  GTECH_XOR2 U166 ( .A(n313), .B(n319), .Z(n318) );
  GTECH_AOI21 U167 ( .A(n320), .B(n321), .C(n322), .Z(n313) );
  GTECH_XOR2 U168 ( .A(n323), .B(n319), .Z(n317) );
  GTECH_XOR2 U169 ( .A(a[2]), .B(b[2]), .Z(n319) );
  GTECH_OAI2N2 U170 ( .A(n324), .B(n325), .C(n326), .D(n325), .Z(sum[1]) );
  GTECH_OAI21 U171 ( .A(cin), .B(n321), .C(n327), .Z(n326) );
  GTECH_AND_NOT U172 ( .A(n320), .B(n322), .Z(n325) );
  GTECH_AOI21 U173 ( .A(n327), .B(cin), .C(n321), .Z(n324) );
  GTECH_OAI22 U174 ( .A(n328), .B(n329), .C(n330), .D(n331), .Z(sum[15]) );
  GTECH_XNOR2 U175 ( .A(n332), .B(n333), .Z(n331) );
  GTECH_XNOR2 U176 ( .A(n333), .B(n334), .Z(n329) );
  GTECH_ADD_ABC U177 ( .A(a[14]), .B(n335), .C(b[14]), .COUT(n334) );
  GTECH_XOR2 U178 ( .A(a[15]), .B(b[15]), .Z(n333) );
  GTECH_OAI22 U179 ( .A(n328), .B(n336), .C(n330), .D(n337), .Z(sum[14]) );
  GTECH_XOR2 U180 ( .A(n338), .B(n339), .Z(n337) );
  GTECH_XOR2 U181 ( .A(n338), .B(n335), .Z(n336) );
  GTECH_OA21 U182 ( .A(n340), .B(n341), .C(n342), .Z(n335) );
  GTECH_XNOR2 U183 ( .A(a[14]), .B(b[14]), .Z(n338) );
  GTECH_OAI22 U184 ( .A(n328), .B(n343), .C(n330), .D(n344), .Z(sum[13]) );
  GTECH_XNOR2 U185 ( .A(n345), .B(n346), .Z(n344) );
  GTECH_XOR2 U186 ( .A(n341), .B(n345), .Z(n343) );
  GTECH_OAI21 U187 ( .A(a[13]), .B(b[13]), .C(n347), .Z(n345) );
  GTECH_NAND2 U188 ( .A(n348), .B(n349), .Z(sum[12]) );
  GTECH_OAI21 U189 ( .A(n341), .B(n346), .C(n328), .Z(n348) );
  GTECH_OAI22 U190 ( .A(n350), .B(n271), .C(n272), .D(n351), .Z(sum[11]) );
  GTECH_XNOR2 U191 ( .A(n352), .B(n353), .Z(n351) );
  GTECH_ADD_ABC U192 ( .A(a[10]), .B(n354), .C(b[10]), .COUT(n353) );
  GTECH_XNOR2 U193 ( .A(n355), .B(n352), .Z(n350) );
  GTECH_XOR2 U194 ( .A(a[11]), .B(b[11]), .Z(n352) );
  GTECH_OAI22 U195 ( .A(n272), .B(n356), .C(n271), .D(n357), .Z(sum[10]) );
  GTECH_XOR2 U196 ( .A(n358), .B(n359), .Z(n357) );
  GTECH_XOR2 U197 ( .A(n358), .B(n354), .Z(n356) );
  GTECH_OA21 U198 ( .A(n360), .B(n274), .C(n361), .Z(n354) );
  GTECH_XNOR2 U199 ( .A(a[10]), .B(b[10]), .Z(n358) );
  GTECH_XOR2 U200 ( .A(cin), .B(n362), .Z(sum[0]) );
  GTECH_OAI21 U201 ( .A(n330), .B(n363), .C(n349), .Z(cout) );
  GTECH_OR3 U202 ( .A(n346), .B(n341), .C(n328), .Z(n349) );
  GTECH_NOT U203 ( .A(n330), .Z(n328) );
  GTECH_AND2 U204 ( .A(b[12]), .B(a[12]), .Z(n341) );
  GTECH_AOI21 U205 ( .A(n332), .B(a[15]), .C(n364), .Z(n363) );
  GTECH_OA21 U206 ( .A(a[15]), .B(n332), .C(b[15]), .Z(n364) );
  GTECH_ADD_ABC U207 ( .A(a[14]), .B(n339), .C(b[14]), .COUT(n332) );
  GTECH_OA21 U208 ( .A(n340), .B(n365), .C(n342), .Z(n339) );
  GTECH_OR2 U209 ( .A(b[13]), .B(a[13]), .Z(n342) );
  GTECH_NOT U210 ( .A(n346), .Z(n365) );
  GTECH_NOR2 U211 ( .A(a[12]), .B(b[12]), .Z(n346) );
  GTECH_NOT U212 ( .A(n347), .Z(n340) );
  GTECH_NAND2 U213 ( .A(b[13]), .B(a[13]), .Z(n347) );
  GTECH_OA21 U214 ( .A(n271), .B(n366), .C(n280), .Z(n330) );
  GTECH_OR_NOT U215 ( .A(n272), .B(n279), .Z(n280) );
  GTECH_AND_NOT U216 ( .A(n277), .B(n274), .Z(n279) );
  GTECH_AND2 U217 ( .A(b[8]), .B(a[8]), .Z(n274) );
  GTECH_OAI21 U218 ( .A(a[11]), .B(n355), .C(n367), .Z(n366) );
  GTECH_NOT U219 ( .A(n368), .Z(n367) );
  GTECH_AOI21 U220 ( .A(n355), .B(a[11]), .C(b[11]), .Z(n368) );
  GTECH_ADD_ABC U221 ( .A(n359), .B(a[10]), .C(b[10]), .COUT(n355) );
  GTECH_OA21 U222 ( .A(n360), .B(n277), .C(n361), .Z(n359) );
  GTECH_OR2 U223 ( .A(b[9]), .B(a[9]), .Z(n361) );
  GTECH_OR2 U224 ( .A(a[8]), .B(b[8]), .Z(n277) );
  GTECH_NOT U225 ( .A(n278), .Z(n360) );
  GTECH_NAND2 U226 ( .A(b[9]), .B(a[9]), .Z(n278) );
  GTECH_NOT U227 ( .A(n272), .Z(n271) );
  GTECH_AOI2N2 U228 ( .A(n306), .B(n284), .C(n369), .D(n284), .Z(n272) );
  GTECH_OA21 U229 ( .A(a[7]), .B(n285), .C(n370), .Z(n369) );
  GTECH_NOT U230 ( .A(n371), .Z(n370) );
  GTECH_AOI21 U231 ( .A(n285), .B(a[7]), .C(b[7]), .Z(n371) );
  GTECH_OAI21 U232 ( .A(n294), .B(n288), .C(n372), .Z(n285) );
  GTECH_OAI21 U233 ( .A(a[6]), .B(n373), .C(b[6]), .Z(n372) );
  GTECH_NOT U234 ( .A(a[6]), .Z(n288) );
  GTECH_NOT U235 ( .A(n373), .Z(n294) );
  GTECH_OAI21 U236 ( .A(n303), .B(n296), .C(n298), .Z(n373) );
  GTECH_NAND2 U237 ( .A(b[5]), .B(a[5]), .Z(n298) );
  GTECH_NOR2 U238 ( .A(a[5]), .B(b[5]), .Z(n296) );
  GTECH_NOR2 U239 ( .A(a[4]), .B(b[4]), .Z(n303) );
  GTECH_AOI2N2 U240 ( .A(n307), .B(n362), .C(n374), .D(n307), .Z(n284) );
  GTECH_AOI21 U241 ( .A(n316), .B(a[3]), .C(n375), .Z(n374) );
  GTECH_OA21 U242 ( .A(a[3]), .B(n316), .C(b[3]), .Z(n375) );
  GTECH_OAI21 U243 ( .A(n323), .B(n312), .C(n376), .Z(n316) );
  GTECH_OAI21 U244 ( .A(a[2]), .B(n377), .C(b[2]), .Z(n376) );
  GTECH_NOT U245 ( .A(n323), .Z(n377) );
  GTECH_NOT U246 ( .A(a[2]), .Z(n312) );
  GTECH_AOI21 U247 ( .A(n327), .B(n320), .C(n322), .Z(n323) );
  GTECH_AND2 U248 ( .A(b[1]), .B(a[1]), .Z(n322) );
  GTECH_OR2 U249 ( .A(b[1]), .B(a[1]), .Z(n320) );
  GTECH_AND_NOT U250 ( .A(n327), .B(n321), .Z(n362) );
  GTECH_AND2 U251 ( .A(b[0]), .B(a[0]), .Z(n321) );
  GTECH_OR2 U252 ( .A(b[0]), .B(a[0]), .Z(n327) );
  GTECH_NOT U253 ( .A(cin), .Z(n307) );
  GTECH_XOR2 U254 ( .A(n304), .B(b[4]), .Z(n306) );
  GTECH_NOT U255 ( .A(a[4]), .Z(n304) );
endmodule

