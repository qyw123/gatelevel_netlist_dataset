
module CRC32 ( crcIn, data, crcOut );
  input [31:0] crcIn;
  input [7:0] data;
  output [31:0] crcOut;
  wire   n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  GTECH_XNOR2 U62 ( .A(crcIn[17]), .B(n30), .Z(crcOut[9]) );
  GTECH_XNOR3 U63 ( .A(crcIn[16]), .B(n31), .C(n32), .Z(crcOut[8]) );
  GTECH_ADD_ABC U64 ( .A(crcIn[15]), .B(n33), .C(n34), .S(crcOut[7]) );
  GTECH_XNOR2 U65 ( .A(crcIn[14]), .B(n35), .Z(crcOut[6]) );
  GTECH_XNOR3 U66 ( .A(crcIn[13]), .B(n36), .C(crcOut[31]), .Z(crcOut[5]) );
  GTECH_ADD_ABC U67 ( .A(crcIn[12]), .B(n33), .C(n37), .S(crcOut[4]) );
  GTECH_ADD_ABC U68 ( .A(crcIn[11]), .B(n38), .C(n39), .S(crcOut[3]) );
  GTECH_ADD_ABC U69 ( .A(crcIn[10]), .B(n40), .C(n41), .S(crcOut[2]) );
  GTECH_XOR2 U70 ( .A(n34), .B(crcOut[30]), .Z(crcOut[29]) );
  GTECH_XOR2 U71 ( .A(n33), .B(n42), .Z(crcOut[28]) );
  GTECH_XOR2 U72 ( .A(n43), .B(n44), .Z(n33) );
  GTECH_XNOR3 U73 ( .A(n35), .B(n45), .C(crcOut[31]), .Z(crcOut[27]) );
  GTECH_XOR2 U74 ( .A(n31), .B(n30), .Z(crcOut[31]) );
  GTECH_ADD_ABC U75 ( .A(n40), .B(n37), .C(crcOut[30]), .S(crcOut[26]) );
  GTECH_XOR2 U76 ( .A(n41), .B(n32), .Z(crcOut[30]) );
  GTECH_XOR2 U77 ( .A(n46), .B(n47), .Z(crcOut[25]) );
  GTECH_NOT U78 ( .A(n41), .Z(n46) );
  GTECH_XOR2 U79 ( .A(n43), .B(n48), .Z(crcOut[24]) );
  GTECH_XNOR2 U80 ( .A(crcIn[31]), .B(n49), .Z(crcOut[23]) );
  GTECH_XNOR2 U81 ( .A(crcIn[30]), .B(n47), .Z(crcOut[22]) );
  GTECH_ADD_ABC U82 ( .A(n44), .B(n34), .C(n37), .S(n47) );
  GTECH_XNOR2 U83 ( .A(crcIn[29]), .B(n48), .Z(crcOut[21]) );
  GTECH_ADD_ABC U84 ( .A(n50), .B(n35), .C(n51), .S(n48) );
  GTECH_XNOR2 U85 ( .A(crcIn[28]), .B(n49), .Z(crcOut[20]) );
  GTECH_XOR2 U86 ( .A(n36), .B(n32), .Z(n49) );
  GTECH_XNOR2 U87 ( .A(n45), .B(n40), .Z(n36) );
  GTECH_ADD_ABC U88 ( .A(crcIn[9]), .B(n52), .C(n45), .S(crcOut[1]) );
  GTECH_XNOR4 U89 ( .A(crcIn[27]), .B(n32), .C(n39), .D(n37), .Z(crcOut[19])
         );
  GTECH_XNOR2 U90 ( .A(n34), .B(n53), .Z(n39) );
  GTECH_XNOR2 U91 ( .A(n44), .B(n50), .Z(n32) );
  GTECH_NOT U92 ( .A(n54), .Z(n44) );
  GTECH_XNOR3 U93 ( .A(crcIn[26]), .B(n55), .C(n56), .Z(crcOut[18]) );
  GTECH_ADD_ABC U94 ( .A(crcIn[25]), .B(n45), .C(n56), .S(crcOut[17]) );
  GTECH_XNOR2 U95 ( .A(n41), .B(n35), .Z(n56) );
  GTECH_NOT U96 ( .A(n42), .Z(n35) );
  GTECH_XOR2 U97 ( .A(n40), .B(n34), .Z(n42) );
  GTECH_ADD_ABC U98 ( .A(crcIn[24]), .B(n37), .C(n57), .S(crcOut[16]) );
  GTECH_XNOR3 U99 ( .A(crcIn[23]), .B(n30), .C(n37), .Z(crcOut[15]) );
  GTECH_XNOR2 U100 ( .A(n38), .B(n45), .Z(n37) );
  GTECH_NOT U101 ( .A(n50), .Z(n30) );
  GTECH_XOR2 U102 ( .A(data[7]), .B(crcIn[7]), .Z(n50) );
  GTECH_ADD_ABC U103 ( .A(crcIn[22]), .B(n31), .C(n55), .S(crcOut[14]) );
  GTECH_XNOR2 U104 ( .A(n51), .B(n54), .Z(n55) );
  GTECH_XOR2 U105 ( .A(data[6]), .B(crcIn[6]), .Z(n54) );
  GTECH_NOT U106 ( .A(n53), .Z(n31) );
  GTECH_ADD_ABC U107 ( .A(crcIn[21]), .B(n34), .C(n41), .S(crcOut[13]) );
  GTECH_XNOR2 U108 ( .A(n43), .B(n53), .Z(n41) );
  GTECH_XOR2 U109 ( .A(data[1]), .B(crcIn[1]), .Z(n53) );
  GTECH_NOT U110 ( .A(n52), .Z(n43) );
  GTECH_XOR2 U111 ( .A(data[5]), .B(crcIn[5]), .Z(n34) );
  GTECH_XOR2 U112 ( .A(crcIn[20]), .B(n57), .Z(crcOut[12]) );
  GTECH_XOR2 U113 ( .A(n40), .B(n52), .Z(n57) );
  GTECH_XOR2 U114 ( .A(data[0]), .B(crcIn[0]), .Z(n52) );
  GTECH_XOR2 U115 ( .A(data[4]), .B(crcIn[4]), .Z(n40) );
  GTECH_XOR2 U116 ( .A(crcIn[19]), .B(n45), .Z(crcOut[11]) );
  GTECH_XOR2 U117 ( .A(data[3]), .B(crcIn[3]), .Z(n45) );
  GTECH_XNOR2 U118 ( .A(crcIn[18]), .B(n38), .Z(crcOut[10]) );
  GTECH_XNOR2 U119 ( .A(crcIn[8]), .B(n38), .Z(crcOut[0]) );
  GTECH_NOT U120 ( .A(n51), .Z(n38) );
  GTECH_XOR2 U121 ( .A(data[2]), .B(crcIn[2]), .Z(n51) );
endmodule

