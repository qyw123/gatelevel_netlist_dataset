
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398;

  GTECH_MUX2 U143 ( .A(n282), .B(n283), .S(n284), .Z(sum[9]) );
  GTECH_OA21 U144 ( .A(n285), .B(n286), .C(n287), .Z(n284) );
  GTECH_OR_NOT U145 ( .A(n288), .B(n289), .Z(n283) );
  GTECH_XOR2 U146 ( .A(b[9]), .B(a[9]), .Z(n282) );
  GTECH_OAI21 U147 ( .A(n290), .B(n291), .C(n292), .Z(sum[8]) );
  GTECH_NOR2 U148 ( .A(n293), .B(n285), .Z(n290) );
  GTECH_MUX2 U149 ( .A(n294), .B(n295), .S(n296), .Z(sum[7]) );
  GTECH_XOR2 U150 ( .A(n297), .B(n298), .Z(n295) );
  GTECH_AND_NOT U151 ( .A(n299), .B(n300), .Z(n298) );
  GTECH_OAI21 U152 ( .A(b[6]), .B(a[6]), .C(n301), .Z(n299) );
  GTECH_XNOR2 U153 ( .A(n297), .B(n302), .Z(n294) );
  GTECH_XNOR2 U154 ( .A(a[7]), .B(b[7]), .Z(n297) );
  GTECH_AO21 U155 ( .A(n303), .B(n300), .C(n304), .Z(sum[6]) );
  GTECH_NOT U156 ( .A(n305), .Z(n304) );
  GTECH_MUX2 U157 ( .A(n306), .B(n307), .S(b[6]), .Z(n305) );
  GTECH_OR_NOT U158 ( .A(n303), .B(n308), .Z(n307) );
  GTECH_XOR2 U159 ( .A(n308), .B(n303), .Z(n306) );
  GTECH_AO21 U160 ( .A(n309), .B(n310), .C(n301), .Z(n303) );
  GTECH_AO21 U161 ( .A(a[4]), .B(n311), .C(n312), .Z(n301) );
  GTECH_AND_NOT U162 ( .A(b[4]), .B(n313), .Z(n311) );
  GTECH_MUX2 U163 ( .A(n314), .B(n315), .S(n316), .Z(sum[5]) );
  GTECH_AND_NOT U164 ( .A(n317), .B(n313), .Z(n316) );
  GTECH_OAI21 U165 ( .A(a[4]), .B(n310), .C(n318), .Z(n315) );
  GTECH_AO21 U166 ( .A(n310), .B(a[4]), .C(b[4]), .Z(n318) );
  GTECH_OAI2N2 U167 ( .A(n319), .B(n296), .C(b[4]), .D(a[4]), .Z(n314) );
  GTECH_XNOR2 U168 ( .A(n320), .B(n296), .Z(sum[4]) );
  GTECH_MUX2 U169 ( .A(n321), .B(n322), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U170 ( .A(n323), .B(n324), .Z(n322) );
  GTECH_XOR2 U171 ( .A(n325), .B(n323), .Z(n321) );
  GTECH_XOR2 U172 ( .A(a[3]), .B(b[3]), .Z(n323) );
  GTECH_OA21 U173 ( .A(a[2]), .B(n326), .C(n327), .Z(n325) );
  GTECH_AO21 U174 ( .A(n326), .B(a[2]), .C(b[2]), .Z(n327) );
  GTECH_MUX2 U175 ( .A(n328), .B(n329), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U176 ( .A(n330), .B(n331), .Z(n329) );
  GTECH_XNOR2 U177 ( .A(n330), .B(n326), .Z(n328) );
  GTECH_AO21 U178 ( .A(n332), .B(n333), .C(n334), .Z(n326) );
  GTECH_XOR2 U179 ( .A(a[2]), .B(n335), .Z(n330) );
  GTECH_MUX2 U180 ( .A(n336), .B(n337), .S(n338), .Z(sum[1]) );
  GTECH_AND_NOT U181 ( .A(n332), .B(n334), .Z(n338) );
  GTECH_OAI21 U182 ( .A(cin), .B(n333), .C(n339), .Z(n337) );
  GTECH_OAI21 U183 ( .A(n340), .B(n341), .C(n342), .Z(n336) );
  GTECH_NOT U184 ( .A(n333), .Z(n342) );
  GTECH_NOT U185 ( .A(cin), .Z(n341) );
  GTECH_MUX2 U186 ( .A(n343), .B(n344), .S(n345), .Z(sum[15]) );
  GTECH_XOR2 U187 ( .A(n346), .B(n347), .Z(n344) );
  GTECH_OA21 U188 ( .A(n348), .B(n349), .C(n350), .Z(n347) );
  GTECH_XNOR2 U189 ( .A(n346), .B(n351), .Z(n343) );
  GTECH_XNOR2 U190 ( .A(a[15]), .B(b[15]), .Z(n346) );
  GTECH_MUX2 U191 ( .A(n352), .B(n353), .S(n345), .Z(sum[14]) );
  GTECH_XNOR2 U192 ( .A(n349), .B(n354), .Z(n353) );
  GTECH_AOI21 U193 ( .A(n355), .B(n356), .C(n357), .Z(n349) );
  GTECH_XNOR2 U194 ( .A(n354), .B(n358), .Z(n352) );
  GTECH_AND_NOT U195 ( .A(n350), .B(n348), .Z(n354) );
  GTECH_MUX2 U196 ( .A(n359), .B(n360), .S(n345), .Z(sum[13]) );
  GTECH_XNOR2 U197 ( .A(n361), .B(n362), .Z(n360) );
  GTECH_XOR2 U198 ( .A(n362), .B(n363), .Z(n359) );
  GTECH_AND_NOT U199 ( .A(n355), .B(n357), .Z(n362) );
  GTECH_OAI21 U200 ( .A(n345), .B(n364), .C(n365), .Z(sum[12]) );
  GTECH_AND2 U201 ( .A(n363), .B(n361), .Z(n364) );
  GTECH_MUX2 U202 ( .A(n366), .B(n367), .S(n291), .Z(sum[11]) );
  GTECH_XOR2 U203 ( .A(n368), .B(n369), .Z(n367) );
  GTECH_AND2 U204 ( .A(n370), .B(n371), .Z(n369) );
  GTECH_OAI21 U205 ( .A(b[10]), .B(a[10]), .C(n372), .Z(n370) );
  GTECH_OA21 U206 ( .A(n285), .B(n288), .C(n289), .Z(n372) );
  GTECH_XNOR2 U207 ( .A(n368), .B(n373), .Z(n366) );
  GTECH_XNOR2 U208 ( .A(a[11]), .B(b[11]), .Z(n368) );
  GTECH_OAI21 U209 ( .A(n374), .B(n371), .C(n375), .Z(sum[10]) );
  GTECH_MUX2 U210 ( .A(n376), .B(n377), .S(b[10]), .Z(n375) );
  GTECH_OR_NOT U211 ( .A(a[10]), .B(n374), .Z(n377) );
  GTECH_XNOR2 U212 ( .A(n378), .B(n374), .Z(n376) );
  GTECH_OA21 U213 ( .A(n291), .B(n379), .C(n380), .Z(n374) );
  GTECH_OAI21 U214 ( .A(n288), .B(n285), .C(n289), .Z(n380) );
  GTECH_XOR2 U215 ( .A(cin), .B(n381), .Z(sum[0]) );
  GTECH_OAI21 U216 ( .A(n345), .B(n382), .C(n365), .Z(cout) );
  GTECH_NAND3 U217 ( .A(n361), .B(n363), .C(n345), .Z(n365) );
  GTECH_NOT U218 ( .A(n356), .Z(n361) );
  GTECH_AND_NOT U219 ( .A(b[12]), .B(n383), .Z(n356) );
  GTECH_AOI21 U220 ( .A(n351), .B(a[15]), .C(n384), .Z(n382) );
  GTECH_OA21 U221 ( .A(a[15]), .B(n351), .C(b[15]), .Z(n384) );
  GTECH_OAI21 U222 ( .A(n358), .B(n348), .C(n350), .Z(n351) );
  GTECH_OR_NOT U223 ( .A(n385), .B(b[14]), .Z(n350) );
  GTECH_AND_NOT U224 ( .A(n385), .B(b[14]), .Z(n348) );
  GTECH_NOT U225 ( .A(a[14]), .Z(n385) );
  GTECH_AOI21 U226 ( .A(n355), .B(n363), .C(n357), .Z(n358) );
  GTECH_AND2 U227 ( .A(a[13]), .B(b[13]), .Z(n357) );
  GTECH_OR_NOT U228 ( .A(b[12]), .B(n383), .Z(n363) );
  GTECH_NOT U229 ( .A(a[12]), .Z(n383) );
  GTECH_NOT U230 ( .A(n386), .Z(n355) );
  GTECH_NOR2 U231 ( .A(a[13]), .B(b[13]), .Z(n386) );
  GTECH_OA21 U232 ( .A(n387), .B(n291), .C(n292), .Z(n345) );
  GTECH_OR3 U233 ( .A(n285), .B(n293), .C(n286), .Z(n292) );
  GTECH_AND2 U234 ( .A(a[8]), .B(b[8]), .Z(n285) );
  GTECH_NOT U235 ( .A(n286), .Z(n291) );
  GTECH_MUX2 U236 ( .A(n388), .B(n320), .S(n296), .Z(n286) );
  GTECH_NOT U237 ( .A(n310), .Z(n296) );
  GTECH_MUX2 U238 ( .A(n381), .B(n389), .S(cin), .Z(n310) );
  GTECH_OA21 U239 ( .A(a[3]), .B(n324), .C(n390), .Z(n389) );
  GTECH_AO21 U240 ( .A(n324), .B(a[3]), .C(b[3]), .Z(n390) );
  GTECH_OAI21 U241 ( .A(n331), .B(n391), .C(n392), .Z(n324) );
  GTECH_AO21 U242 ( .A(n391), .B(n331), .C(n335), .Z(n392) );
  GTECH_NOT U243 ( .A(b[2]), .Z(n335) );
  GTECH_NOT U244 ( .A(a[2]), .Z(n391) );
  GTECH_AOI21 U245 ( .A(n332), .B(n339), .C(n334), .Z(n331) );
  GTECH_AND2 U246 ( .A(a[1]), .B(b[1]), .Z(n334) );
  GTECH_NOT U247 ( .A(n393), .Z(n332) );
  GTECH_NOR2 U248 ( .A(a[1]), .B(b[1]), .Z(n393) );
  GTECH_AND_NOT U249 ( .A(n339), .B(n333), .Z(n381) );
  GTECH_AND2 U250 ( .A(a[0]), .B(b[0]), .Z(n333) );
  GTECH_NOT U251 ( .A(n340), .Z(n339) );
  GTECH_NOR2 U252 ( .A(a[0]), .B(b[0]), .Z(n340) );
  GTECH_XOR2 U253 ( .A(a[4]), .B(b[4]), .Z(n320) );
  GTECH_OA21 U254 ( .A(a[7]), .B(n302), .C(n394), .Z(n388) );
  GTECH_AO21 U255 ( .A(n302), .B(a[7]), .C(b[7]), .Z(n394) );
  GTECH_AO21 U256 ( .A(n309), .B(n395), .C(n300), .Z(n302) );
  GTECH_AND_NOT U257 ( .A(b[6]), .B(n308), .Z(n300) );
  GTECH_OR_NOT U258 ( .A(b[6]), .B(n308), .Z(n395) );
  GTECH_NOT U259 ( .A(a[6]), .Z(n308) );
  GTECH_OAI21 U260 ( .A(n313), .B(n319), .C(n317), .Z(n309) );
  GTECH_NOT U261 ( .A(n312), .Z(n317) );
  GTECH_AND2 U262 ( .A(a[5]), .B(b[5]), .Z(n312) );
  GTECH_NOR2 U263 ( .A(a[4]), .B(b[4]), .Z(n319) );
  GTECH_NOR2 U264 ( .A(a[5]), .B(b[5]), .Z(n313) );
  GTECH_AOI21 U265 ( .A(n373), .B(a[11]), .C(n396), .Z(n387) );
  GTECH_OA21 U266 ( .A(a[11]), .B(n373), .C(b[11]), .Z(n396) );
  GTECH_OAI21 U267 ( .A(n397), .B(n379), .C(n371), .Z(n373) );
  GTECH_OR_NOT U268 ( .A(n378), .B(b[10]), .Z(n371) );
  GTECH_NOT U269 ( .A(a[10]), .Z(n378) );
  GTECH_OAI21 U270 ( .A(n288), .B(n287), .C(n289), .Z(n379) );
  GTECH_NOT U271 ( .A(n398), .Z(n289) );
  GTECH_NOR2 U272 ( .A(a[9]), .B(b[9]), .Z(n398) );
  GTECH_NOT U273 ( .A(n293), .Z(n287) );
  GTECH_NOR2 U274 ( .A(a[8]), .B(b[8]), .Z(n293) );
  GTECH_AND2 U275 ( .A(a[9]), .B(b[9]), .Z(n288) );
  GTECH_NOR2 U276 ( .A(a[10]), .B(b[10]), .Z(n397) );
endmodule

