
module frequency_counter ( clk, reset, signal, period, period_load, segments, 
        digit, dbg_state, dbg_clk_count, dbg_edge_count );
  input [11:0] period;
  output [6:0] segments;
  output [1:0] dbg_state;
  output [2:0] dbg_clk_count;
  output [2:0] dbg_edge_count;
  input clk, reset, signal, period_load;
  output digit;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21,
         update_digits, N62, N112, N114, N116, N118, N120, N122, N124, N126,
         N128, N130, N132, N133, N134, N136, N138, N140, N142, N144, N146,
         N147, N148, N150, N151, N152, N154, N156, N158, N159, N160, N162,
         N164, N166, N167, N168, N169, N170, edge_detect0_q2, edge_detect0_q1,
         edge_detect0_q0, seven_segment0_N22, seven_segment0_N20,
         seven_segment0_N18, seven_segment0_N16, seven_segment0_N14,
         seven_segment0_N12, seven_segment0_N10, seven_segment0_N9,
         seven_segment0_N8, seven_segment0_N6, n13, n14, n15, n16, n20, n22,
         n27, n28, n29, n31, n32, n33, n78, n156, n159, sub_85_carry_2_, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n175, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353;
  wire   [8:0] clk_counter;
  wire   [3:0] edge_counter;
  wire   [11:0] update_period;
  wire   [3:0] ten_count;
  wire   [3:0] unit_count;
  wire   [0:3] seven_segment0_unit_count_reg;
  wire   [0:3] seven_segment0_ten_count_reg;

  GTECH_FJK1S update_period_reg_11_ ( .J(n78), .K(n78), .TI(N21), .TE(N20), 
        .CP(clk), .Q(update_period[11]) );
  GTECH_FJK1S update_period_reg_10_ ( .J(n78), .K(n78), .TI(N19), .TE(N20), 
        .CP(clk), .Q(update_period[10]) );
  GTECH_FJK1S update_period_reg_9_ ( .J(n78), .K(n78), .TI(N18), .TE(N20), 
        .CP(clk), .Q(update_period[9]) );
  GTECH_FJK1S update_period_reg_8_ ( .J(n78), .K(n78), .TI(N17), .TE(N20), 
        .CP(clk), .Q(update_period[8]) );
  GTECH_FJK1S update_period_reg_7_ ( .J(n78), .K(n78), .TI(N16), .TE(N20), 
        .CP(clk), .Q(update_period[7]) );
  GTECH_FJK1S update_period_reg_6_ ( .J(n78), .K(n78), .TI(N15), .TE(N20), 
        .CP(clk), .Q(update_period[6]) );
  GTECH_FJK1S update_period_reg_5_ ( .J(n78), .K(n78), .TI(N14), .TE(N20), 
        .CP(clk), .Q(update_period[5]) );
  GTECH_FJK1S update_period_reg_4_ ( .J(n78), .K(n78), .TI(N13), .TE(N20), 
        .CP(clk), .Q(update_period[4]) );
  GTECH_FJK1S update_period_reg_3_ ( .J(n78), .K(n78), .TI(N12), .TE(N20), 
        .CP(clk), .Q(update_period[3]) );
  GTECH_FJK1S update_period_reg_2_ ( .J(n78), .K(n78), .TI(N11), .TE(N20), 
        .CP(clk), .Q(update_period[2]) );
  GTECH_FJK1S update_period_reg_1_ ( .J(n78), .K(n78), .TI(N10), .TE(N20), 
        .CP(clk), .Q(update_period[1]), .QN(n175) );
  GTECH_FJK1S update_period_reg_0_ ( .J(n78), .K(n78), .TI(N9), .TE(N20), .CP(
        clk), .Q(update_period[0]) );
  GTECH_FD1 edge_detect0_q0_reg ( .D(signal), .CP(clk), .Q(edge_detect0_q0) );
  GTECH_FD1 edge_detect0_q1_reg ( .D(edge_detect0_q0), .CP(clk), .Q(
        edge_detect0_q1) );
  GTECH_FD1 edge_detect0_q2_reg ( .D(edge_detect0_q1), .CP(clk), .Q(
        edge_detect0_q2), .QN(n13) );
  GTECH_FJK1S edge_counter_reg_5_ ( .J(n78), .K(n78), .TI(N146), .TE(N147), 
        .CP(clk), .Q(dbg_edge_count[1]), .QN(n173) );
  GTECH_FJK1S edge_counter_reg_6_ ( .J(n78), .K(n78), .TI(N148), .TE(N147), 
        .CP(clk), .Q(dbg_edge_count[2]), .QN(n172) );
  GTECH_FJK1S state_reg_0_ ( .J(n78), .K(n78), .TI(N150), .TE(N151), .CP(clk), 
        .Q(dbg_state[0]), .QN(n14) );
  GTECH_FJK1S state_reg_1_ ( .J(n78), .K(n78), .TI(N152), .TE(N151), .CP(clk), 
        .Q(dbg_state[1]), .QN(n159) );
  GTECH_FJK1S update_digits_reg ( .J(n78), .K(n78), .TI(N170), .TE(N169), .CP(
        clk), .Q(update_digits), .QN(n15) );
  GTECH_FJK1S clk_counter_reg_10_ ( .J(n78), .K(n78), .TI(N132), .TE(N133), 
        .CP(clk), .Q(dbg_clk_count[1]), .QN(n171) );
  GTECH_FJK1S clk_counter_reg_0_ ( .J(n78), .K(n78), .TI(N112), .TE(N133), 
        .CP(clk), .Q(clk_counter[0]), .QN(n170) );
  GTECH_FJK1S clk_counter_reg_1_ ( .J(n78), .K(n78), .TI(N114), .TE(N133), 
        .CP(clk), .Q(clk_counter[1]), .QN(n169) );
  GTECH_FJK1S clk_counter_reg_2_ ( .J(n78), .K(n78), .TI(N116), .TE(N133), 
        .CP(clk), .Q(clk_counter[2]), .QN(n168) );
  GTECH_FJK1S clk_counter_reg_3_ ( .J(n78), .K(n78), .TI(N118), .TE(N133), 
        .CP(clk), .Q(clk_counter[3]), .QN(n167) );
  GTECH_FJK1S clk_counter_reg_4_ ( .J(n78), .K(n78), .TI(N120), .TE(N133), 
        .CP(clk), .Q(clk_counter[4]), .QN(n166) );
  GTECH_FJK1S clk_counter_reg_5_ ( .J(n78), .K(n78), .TI(N122), .TE(N133), 
        .CP(clk), .Q(clk_counter[5]), .QN(n165) );
  GTECH_FJK1S clk_counter_reg_6_ ( .J(n78), .K(n78), .TI(N124), .TE(N133), 
        .CP(clk), .Q(clk_counter[6]), .QN(n164) );
  GTECH_FJK1S clk_counter_reg_7_ ( .J(n78), .K(n78), .TI(N126), .TE(N133), 
        .CP(clk), .Q(clk_counter[7]), .QN(n163) );
  GTECH_FJK1S clk_counter_reg_8_ ( .J(n78), .K(n78), .TI(N128), .TE(N133), 
        .CP(clk), .Q(clk_counter[8]), .QN(n162) );
  GTECH_FJK1S clk_counter_reg_9_ ( .J(n78), .K(n78), .TI(N130), .TE(N133), 
        .CP(clk), .Q(dbg_clk_count[0]), .QN(n161) );
  GTECH_FJK1S clk_counter_reg_11_ ( .J(n78), .K(n78), .TI(N134), .TE(N133), 
        .CP(clk), .Q(dbg_clk_count[2]), .QN(n160) );
  GTECH_FJK1S edge_counter_reg_4_ ( .J(n78), .K(n78), .TI(N144), .TE(N147), 
        .CP(clk), .Q(dbg_edge_count[0]), .QN(n186) );
  GTECH_FJK1S edge_counter_reg_0_ ( .J(n78), .K(n78), .TI(N136), .TE(N147), 
        .CP(clk), .Q(N62), .QN(n16) );
  GTECH_FJK1S unit_count_reg_0_ ( .J(n78), .K(n78), .TI(N162), .TE(N167), .CP(
        clk), .Q(unit_count[0]) );
  GTECH_FJK1S edge_counter_reg_1_ ( .J(n78), .K(n78), .TI(N138), .TE(N147), 
        .CP(clk), .Q(sub_85_carry_2_) );
  GTECH_FJK1S unit_count_reg_1_ ( .J(n78), .K(n78), .TI(N164), .TE(N167), .CP(
        clk), .Q(unit_count[1]) );
  GTECH_FJK1S edge_counter_reg_2_ ( .J(n78), .K(n78), .TI(N140), .TE(N147), 
        .CP(clk), .Q(edge_counter[2]), .QN(n20) );
  GTECH_FJK1S unit_count_reg_2_ ( .J(n78), .K(n78), .TI(N166), .TE(N167), .CP(
        clk), .Q(unit_count[2]) );
  GTECH_FJK1S edge_counter_reg_3_ ( .J(n78), .K(n78), .TI(N142), .TE(N147), 
        .CP(clk), .Q(edge_counter[3]), .QN(n22) );
  GTECH_FJK1S unit_count_reg_3_ ( .J(n78), .K(n78), .TI(N168), .TE(N167), .CP(
        clk), .Q(unit_count[3]) );
  GTECH_FJK1S ten_count_reg_0_ ( .J(n78), .K(n78), .TI(N154), .TE(N159), .CP(
        clk), .Q(ten_count[0]) );
  GTECH_FJK1S ten_count_reg_1_ ( .J(n78), .K(n78), .TI(N156), .TE(N159), .CP(
        clk), .Q(ten_count[1]) );
  GTECH_FJK1S ten_count_reg_2_ ( .J(n78), .K(n78), .TI(N158), .TE(N159), .CP(
        clk), .Q(ten_count[2]) );
  GTECH_FJK1S ten_count_reg_3_ ( .J(n78), .K(n78), .TI(N160), .TE(N159), .CP(
        clk), .Q(ten_count[3]) );
  GTECH_FJK1S seven_segment0_unit_count_reg_reg_0_ ( .J(n78), .K(n78), .TI(
        seven_segment0_N16), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_unit_count_reg[0]) );
  GTECH_FJK1S seven_segment0_unit_count_reg_reg_1_ ( .J(n78), .K(n78), .TI(
        seven_segment0_N18), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_unit_count_reg[1]), .QN(n27) );
  GTECH_FJK1S seven_segment0_unit_count_reg_reg_2_ ( .J(n78), .K(n78), .TI(
        seven_segment0_N20), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_unit_count_reg[2]), .QN(n28) );
  GTECH_FJK1S seven_segment0_unit_count_reg_reg_3_ ( .J(n78), .K(n78), .TI(
        seven_segment0_N22), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_unit_count_reg[3]), .QN(n29) );
  GTECH_FJK1S seven_segment0_ten_count_reg_reg_0_ ( .J(n78), .K(n78), .TI(
        seven_segment0_N8), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_ten_count_reg[0]) );
  GTECH_FJK1S seven_segment0_ten_count_reg_reg_1_ ( .J(n78), .K(n78), .TI(
        seven_segment0_N10), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_ten_count_reg[1]), .QN(n31) );
  GTECH_FJK1S seven_segment0_ten_count_reg_reg_2_ ( .J(n78), .K(n78), .TI(
        seven_segment0_N12), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_ten_count_reg[2]), .QN(n32) );
  GTECH_FJK1S seven_segment0_ten_count_reg_reg_3_ ( .J(n78), .K(n78), .TI(
        seven_segment0_N14), .TE(seven_segment0_N9), .CP(clk), .Q(
        seven_segment0_ten_count_reg[3]), .QN(n33) );
  GTECH_FD1 seven_segment0_digit_reg ( .D(seven_segment0_N6), .CP(clk), .Q(
        digit), .QN(n156) );
  GTECH_ZERO U168 ( .Z(n78) );
  GTECH_NAND2 U169 ( .A(n15), .B(n187), .Z(seven_segment0_N9) );
  GTECH_AND2 U170 ( .A(ten_count[0]), .B(n187), .Z(seven_segment0_N8) );
  GTECH_AND2 U171 ( .A(n156), .B(n187), .Z(seven_segment0_N6) );
  GTECH_AND2 U172 ( .A(unit_count[3]), .B(n187), .Z(seven_segment0_N22) );
  GTECH_AND2 U173 ( .A(unit_count[2]), .B(n187), .Z(seven_segment0_N20) );
  GTECH_AND2 U174 ( .A(unit_count[1]), .B(n187), .Z(seven_segment0_N18) );
  GTECH_AND2 U175 ( .A(unit_count[0]), .B(n187), .Z(seven_segment0_N16) );
  GTECH_AND2 U176 ( .A(ten_count[3]), .B(n187), .Z(seven_segment0_N14) );
  GTECH_AND2 U177 ( .A(ten_count[2]), .B(n187), .Z(seven_segment0_N12) );
  GTECH_AND2 U178 ( .A(ten_count[1]), .B(n187), .Z(seven_segment0_N10) );
  GTECH_NAND2 U179 ( .A(n188), .B(n189), .Z(segments[6]) );
  GTECH_OAI21 U180 ( .A(n190), .B(n191), .C(n192), .Z(segments[3]) );
  GTECH_AND_NOT U181 ( .A(n193), .B(segments[4]), .Z(n192) );
  GTECH_OAI21 U182 ( .A(n194), .B(n191), .C(n195), .Z(segments[4]) );
  GTECH_NAND2 U183 ( .A(n196), .B(n197), .Z(segments[2]) );
  GTECH_NOT U184 ( .A(segments[5]), .Z(n197) );
  GTECH_NAND2 U185 ( .A(n198), .B(n189), .Z(segments[5]) );
  GTECH_AND2 U186 ( .A(n193), .B(n199), .Z(n189) );
  GTECH_OR3 U187 ( .A(n194), .B(n200), .C(n201), .Z(n199) );
  GTECH_OA21 U188 ( .A(n202), .B(n203), .C(n195), .Z(n198) );
  GTECH_NOT U189 ( .A(n204), .Z(n196) );
  GTECH_OR3 U190 ( .A(n205), .B(n206), .C(n204), .Z(segments[1]) );
  GTECH_NAND2 U191 ( .A(n207), .B(n203), .Z(n204) );
  GTECH_AND3 U192 ( .A(n202), .B(n208), .C(n209), .Z(n205) );
  GTECH_NAND4 U193 ( .A(n188), .B(n207), .C(n195), .D(n193), .Z(segments[0])
         );
  GTECH_NAND4 U194 ( .A(n209), .B(n194), .C(n202), .D(n190), .Z(n193) );
  GTECH_NAND2 U195 ( .A(n210), .B(n208), .Z(n195) );
  GTECH_NOT U196 ( .A(n203), .Z(n210) );
  GTECH_NAND2 U197 ( .A(n194), .B(n211), .Z(n207) );
  GTECH_NOT U198 ( .A(n191), .Z(n211) );
  GTECH_NOT U199 ( .A(n208), .Z(n194) );
  GTECH_OAI22 U200 ( .A(seven_segment0_ten_count_reg[0]), .B(n156), .C(
        seven_segment0_unit_count_reg[0]), .D(n212), .Z(n208) );
  GTECH_NOT U201 ( .A(n206), .Z(n188) );
  GTECH_OAI22 U202 ( .A(n202), .B(n203), .C(n190), .D(n191), .Z(n206) );
  GTECH_NAND2 U203 ( .A(n202), .B(n213), .Z(n191) );
  GTECH_NAND2 U204 ( .A(n209), .B(n201), .Z(n203) );
  GTECH_NOT U205 ( .A(n190), .Z(n201) );
  GTECH_OAI22 U206 ( .A(n212), .B(n28), .C(n156), .D(n32), .Z(n190) );
  GTECH_NOT U207 ( .A(n213), .Z(n209) );
  GTECH_OAI22 U208 ( .A(n212), .B(n27), .C(n156), .D(n31), .Z(n213) );
  GTECH_NOT U209 ( .A(n200), .Z(n202) );
  GTECH_OAI22 U210 ( .A(n212), .B(n29), .C(n156), .D(n33), .Z(n200) );
  GTECH_NOT U211 ( .A(n156), .Z(n212) );
  GTECH_AO21 U212 ( .A(period[0]), .B(n214), .C(reset), .Z(N9) );
  GTECH_AND2 U213 ( .A(period[11]), .B(n214), .Z(N21) );
  GTECH_NAND2 U214 ( .A(n187), .B(n215), .Z(N20) );
  GTECH_AO21 U215 ( .A(period[10]), .B(n214), .C(reset), .Z(N19) );
  GTECH_AND2 U216 ( .A(period[9]), .B(n214), .Z(N18) );
  GTECH_AND2 U217 ( .A(period[8]), .B(n214), .Z(N17) );
  GTECH_AND2 U218 ( .A(N170), .B(n216), .Z(N168) );
  GTECH_NAND2 U219 ( .A(n217), .B(n218), .Z(N167) );
  GTECH_AND2 U220 ( .A(N170), .B(n219), .Z(N166) );
  GTECH_NOT U221 ( .A(n20), .Z(n219) );
  GTECH_AND2 U222 ( .A(sub_85_carry_2_), .B(N170), .Z(N164) );
  GTECH_AND2 U223 ( .A(N170), .B(n220), .Z(N162) );
  GTECH_NOT U224 ( .A(n221), .Z(N170) );
  GTECH_NAND2 U225 ( .A(n222), .B(n187), .Z(n221) );
  GTECH_OAI22 U226 ( .A(n223), .B(n224), .C(n225), .D(n226), .Z(N160) );
  GTECH_OAI21 U227 ( .A(ten_count[3]), .B(ten_count[2]), .C(n227), .Z(n226) );
  GTECH_OAI21 U228 ( .A(ten_count[3]), .B(n228), .C(ten_count[2]), .Z(n227) );
  GTECH_NOT U229 ( .A(ten_count[3]), .Z(n223) );
  GTECH_AO21 U230 ( .A(period[7]), .B(n214), .C(reset), .Z(N16) );
  GTECH_OAI21 U231 ( .A(n229), .B(n230), .C(n231), .Z(N159) );
  GTECH_NOT U232 ( .A(n232), .Z(n231) );
  GTECH_OAI21 U233 ( .A(n233), .B(n224), .C(n234), .Z(N158) );
  GTECH_OR3 U234 ( .A(n228), .B(n225), .C(ten_count[2]), .Z(n234) );
  GTECH_NAND2 U235 ( .A(N152), .B(n228), .Z(n224) );
  GTECH_NAND2 U236 ( .A(ten_count[1]), .B(ten_count[0]), .Z(n228) );
  GTECH_NOT U237 ( .A(ten_count[2]), .Z(n233) );
  GTECH_OAI21 U238 ( .A(n235), .B(n236), .C(n237), .Z(N156) );
  GTECH_OR3 U239 ( .A(n238), .B(n225), .C(ten_count[1]), .Z(n237) );
  GTECH_NOT U240 ( .A(ten_count[1]), .Z(n235) );
  GTECH_NOT U241 ( .A(n236), .Z(N154) );
  GTECH_NAND2 U242 ( .A(N152), .B(n238), .Z(n236) );
  GTECH_NOT U243 ( .A(ten_count[0]), .Z(n238) );
  GTECH_NAND2 U244 ( .A(n239), .B(n159), .Z(N151) );
  GTECH_OA21 U245 ( .A(n14), .B(n240), .C(n217), .Z(n239) );
  GTECH_NOT U246 ( .A(n241), .Z(n217) );
  GTECH_OAI21 U247 ( .A(n242), .B(n229), .C(n187), .Z(n241) );
  GTECH_AND2 U248 ( .A(period[6]), .B(n214), .Z(N15) );
  GTECH_OAI21 U249 ( .A(n225), .B(n240), .C(n243), .Z(N148) );
  GTECH_AND2 U250 ( .A(n244), .B(n245), .Z(n243) );
  GTECH_NAND4 U251 ( .A(n246), .B(N150), .C(n247), .D(n172), .Z(n245) );
  GTECH_AO21 U252 ( .A(n248), .B(n249), .C(n172), .Z(n244) );
  GTECH_OA22 U253 ( .A(n250), .B(n246), .C(n225), .D(n173), .Z(n248) );
  GTECH_OR3 U254 ( .A(n222), .B(n251), .C(n232), .Z(N147) );
  GTECH_NAND2 U255 ( .A(n187), .B(n252), .Z(n232) );
  GTECH_OR3 U256 ( .A(n14), .B(n253), .C(n254), .Z(n252) );
  GTECH_NOT U257 ( .A(n240), .Z(n253) );
  GTECH_NAND4 U258 ( .A(n186), .B(n173), .C(n172), .D(n255), .Z(n240) );
  GTECH_AND3 U259 ( .A(n14), .B(edge_detect0_q1), .C(n13), .Z(n251) );
  GTECH_NOT U260 ( .A(n218), .Z(n222) );
  GTECH_NAND2 U261 ( .A(n14), .B(n254), .Z(n218) );
  GTECH_NOT U262 ( .A(n159), .Z(n254) );
  GTECH_OAI22 U263 ( .A(n256), .B(n246), .C(n173), .D(n249), .Z(N146) );
  GTECH_OA21 U264 ( .A(n247), .B(n250), .C(n257), .Z(n249) );
  GTECH_OAI21 U265 ( .A(n258), .B(n259), .C(N152), .Z(n257) );
  GTECH_NOT U266 ( .A(n260), .Z(n247) );
  GTECH_NOT U267 ( .A(n173), .Z(n246) );
  GTECH_OA21 U268 ( .A(n260), .B(n250), .C(n261), .Z(n256) );
  GTECH_OR3 U269 ( .A(n186), .B(n22), .C(n262), .Z(n260) );
  GTECH_NAND2 U270 ( .A(n263), .B(n261), .Z(N144) );
  GTECH_OR3 U271 ( .A(n258), .B(n225), .C(n259), .Z(n261) );
  GTECH_NOT U272 ( .A(n186), .Z(n259) );
  GTECH_NOT U273 ( .A(n255), .Z(n258) );
  GTECH_OA21 U274 ( .A(n186), .B(n264), .C(n265), .Z(n263) );
  GTECH_NAND4 U275 ( .A(n266), .B(n216), .C(N150), .D(n186), .Z(n265) );
  GTECH_NOT U276 ( .A(n262), .Z(n266) );
  GTECH_OA21 U277 ( .A(n225), .B(n255), .C(n267), .Z(n264) );
  GTECH_OAI21 U278 ( .A(n22), .B(n262), .C(N150), .Z(n267) );
  GTECH_NAND2 U279 ( .A(n268), .B(n216), .Z(n255) );
  GTECH_NOT U280 ( .A(n269), .Z(N142) );
  GTECH_AOI222 U281 ( .A(n270), .B(N150), .C(n271), .D(n216), .E(n272), .F(n22), .Z(n269) );
  GTECH_AND2 U282 ( .A(N152), .B(n268), .Z(n272) );
  GTECH_NOT U283 ( .A(n22), .Z(n216) );
  GTECH_XOR2 U284 ( .A(n262), .B(n22), .Z(n270) );
  GTECH_OR3 U285 ( .A(n20), .B(n16), .C(n273), .Z(n262) );
  GTECH_OR3 U286 ( .A(n274), .B(n271), .C(n275), .Z(N140) );
  GTECH_AOI21 U287 ( .A(n276), .B(n277), .C(n20), .Z(n275) );
  GTECH_OA22 U288 ( .A(sub_85_carry_2_), .B(n250), .C(n273), .D(n225), .Z(n277) );
  GTECH_NOT U289 ( .A(n278), .Z(n271) );
  GTECH_NAND2 U290 ( .A(n279), .B(N152), .Z(n278) );
  GTECH_NOT U291 ( .A(n225), .Z(N152) );
  GTECH_NOT U292 ( .A(n268), .Z(n279) );
  GTECH_NAND2 U293 ( .A(n20), .B(n273), .Z(n268) );
  GTECH_AND4 U294 ( .A(sub_85_carry_2_), .B(n220), .C(N150), .D(n20), .Z(n274)
         );
  GTECH_NOT U295 ( .A(n16), .Z(n220) );
  GTECH_AO21 U296 ( .A(period[5]), .B(n214), .C(reset), .Z(N14) );
  GTECH_OAI22 U297 ( .A(sub_85_carry_2_), .B(n280), .C(n273), .D(n276), .Z(
        N138) );
  GTECH_NOT U298 ( .A(sub_85_carry_2_), .Z(n273) );
  GTECH_OA21 U299 ( .A(n16), .B(n250), .C(n225), .Z(n280) );
  GTECH_OAI21 U300 ( .A(n16), .B(n225), .C(n276), .Z(N136) );
  GTECH_NAND2 U301 ( .A(n16), .B(N150), .Z(n276) );
  GTECH_NOT U302 ( .A(n250), .Z(N150) );
  GTECH_NAND2 U303 ( .A(n281), .B(n187), .Z(n250) );
  GTECH_NOT U304 ( .A(n230), .Z(n281) );
  GTECH_NAND2 U305 ( .A(n159), .B(n282), .Z(n225) );
  GTECH_NOT U306 ( .A(N169), .Z(n282) );
  GTECH_NAND2 U307 ( .A(n187), .B(n242), .Z(N169) );
  GTECH_NOT U308 ( .A(n14), .Z(n242) );
  GTECH_AND2 U309 ( .A(n283), .B(n284), .Z(N134) );
  GTECH_OAI21 U310 ( .A(n171), .B(n285), .C(n160), .Z(n284) );
  GTECH_NAND2 U311 ( .A(n187), .B(n230), .Z(N133) );
  GTECH_NAND2 U312 ( .A(n159), .B(n14), .Z(n230) );
  GTECH_AND2 U313 ( .A(n286), .B(n283), .Z(N132) );
  GTECH_XOR2 U314 ( .A(n285), .B(n171), .Z(n286) );
  GTECH_NAND2 U315 ( .A(n287), .B(n288), .Z(n285) );
  GTECH_NOT U316 ( .A(n161), .Z(n288) );
  GTECH_NOT U317 ( .A(n289), .Z(n287) );
  GTECH_AND2 U318 ( .A(n290), .B(n283), .Z(N130) );
  GTECH_XOR2 U319 ( .A(n289), .B(n161), .Z(n290) );
  GTECH_NAND2 U320 ( .A(n291), .B(n292), .Z(n289) );
  GTECH_NOT U321 ( .A(n162), .Z(n292) );
  GTECH_NOT U322 ( .A(n293), .Z(n291) );
  GTECH_AND2 U323 ( .A(period[4]), .B(n214), .Z(N13) );
  GTECH_AND2 U324 ( .A(n294), .B(n283), .Z(N128) );
  GTECH_XOR2 U325 ( .A(n293), .B(n162), .Z(n294) );
  GTECH_NAND2 U326 ( .A(n295), .B(n296), .Z(n293) );
  GTECH_NOT U327 ( .A(n297), .Z(n295) );
  GTECH_AND2 U328 ( .A(n298), .B(n283), .Z(N126) );
  GTECH_XOR2 U329 ( .A(n297), .B(n163), .Z(n298) );
  GTECH_NAND2 U330 ( .A(n299), .B(n300), .Z(n297) );
  GTECH_NOT U331 ( .A(n164), .Z(n300) );
  GTECH_NOT U332 ( .A(n301), .Z(n299) );
  GTECH_AND2 U333 ( .A(n302), .B(n283), .Z(N124) );
  GTECH_XOR2 U334 ( .A(n301), .B(n164), .Z(n302) );
  GTECH_NAND2 U335 ( .A(n303), .B(n304), .Z(n301) );
  GTECH_NOT U336 ( .A(n165), .Z(n304) );
  GTECH_NOT U337 ( .A(n305), .Z(n303) );
  GTECH_AND2 U338 ( .A(n306), .B(n283), .Z(N122) );
  GTECH_XOR2 U339 ( .A(n305), .B(n165), .Z(n306) );
  GTECH_NAND2 U340 ( .A(n307), .B(n308), .Z(n305) );
  GTECH_NOT U341 ( .A(n166), .Z(n308) );
  GTECH_NOT U342 ( .A(n309), .Z(n307) );
  GTECH_AND2 U343 ( .A(n310), .B(n283), .Z(N120) );
  GTECH_XOR2 U344 ( .A(n309), .B(n166), .Z(n310) );
  GTECH_NAND2 U345 ( .A(n311), .B(n312), .Z(n309) );
  GTECH_NOT U346 ( .A(n313), .Z(n311) );
  GTECH_AO21 U347 ( .A(period[3]), .B(n214), .C(reset), .Z(N12) );
  GTECH_AND2 U348 ( .A(n314), .B(n283), .Z(N118) );
  GTECH_XOR2 U349 ( .A(n313), .B(n167), .Z(n314) );
  GTECH_OR3 U350 ( .A(n170), .B(n169), .C(n168), .Z(n313) );
  GTECH_OAI22 U351 ( .A(n168), .B(n315), .C(n316), .D(n317), .Z(N116) );
  GTECH_OAI21 U352 ( .A(n169), .B(n168), .C(n318), .Z(n317) );
  GTECH_OAI21 U353 ( .A(n170), .B(n169), .C(n168), .Z(n318) );
  GTECH_OAI21 U354 ( .A(n169), .B(n315), .C(n319), .Z(N114) );
  GTECH_OR3 U355 ( .A(n170), .B(n316), .C(n320), .Z(n319) );
  GTECH_NOT U356 ( .A(n315), .Z(N112) );
  GTECH_NAND2 U357 ( .A(n283), .B(n170), .Z(n315) );
  GTECH_NOT U358 ( .A(n316), .Z(n283) );
  GTECH_NAND2 U359 ( .A(n229), .B(n187), .Z(n316) );
  GTECH_NOT U360 ( .A(n321), .Z(n229) );
  GTECH_AOI222 U361 ( .A(n322), .B(n323), .C(update_period[11]), .D(n160), .E(
        n324), .F(n325), .Z(n321) );
  GTECH_OAI2N2 U362 ( .A(n326), .B(n327), .C(n328), .D(n329), .Z(n324) );
  GTECH_AO22 U363 ( .A(update_period[8]), .B(n330), .C(n161), .D(
        update_period[9]), .Z(n329) );
  GTECH_OA21 U364 ( .A(n161), .B(update_period[9]), .C(n162), .Z(n330) );
  GTECH_OA21 U365 ( .A(n331), .B(n332), .C(n333), .Z(n323) );
  GTECH_AND2 U366 ( .A(n328), .B(n325), .Z(n333) );
  GTECH_NAND2 U367 ( .A(n334), .B(n335), .Z(n325) );
  GTECH_NOT U368 ( .A(update_period[11]), .Z(n335) );
  GTECH_NOT U369 ( .A(n160), .Z(n334) );
  GTECH_NAND2 U370 ( .A(n327), .B(n326), .Z(n328) );
  GTECH_NOT U371 ( .A(n171), .Z(n326) );
  GTECH_NOT U372 ( .A(update_period[10]), .Z(n327) );
  GTECH_OAI2N2 U373 ( .A(n296), .B(n336), .C(n337), .D(n338), .Z(n332) );
  GTECH_AND2 U374 ( .A(update_period[6]), .B(n164), .Z(n337) );
  GTECH_OAI2N2 U375 ( .A(n339), .B(n340), .C(n341), .D(n342), .Z(n331) );
  GTECH_ADD_ABC U376 ( .A(n343), .B(n165), .C(update_period[5]), .COUT(n342)
         );
  GTECH_AND2 U377 ( .A(update_period[4]), .B(n166), .Z(n343) );
  GTECH_OAI21 U378 ( .A(update_period[4]), .B(n166), .C(n341), .Z(n340) );
  GTECH_NOT U379 ( .A(n344), .Z(n341) );
  GTECH_OAI21 U380 ( .A(update_period[6]), .B(n164), .C(n338), .Z(n344) );
  GTECH_NAND2 U381 ( .A(n336), .B(n296), .Z(n338) );
  GTECH_NOT U382 ( .A(n163), .Z(n296) );
  GTECH_NOT U383 ( .A(update_period[7]), .Z(n336) );
  GTECH_OAI22 U384 ( .A(update_period[5]), .B(n165), .C(n345), .D(n346), .Z(
        n339) );
  GTECH_OAI2N2 U385 ( .A(n312), .B(n347), .C(n348), .D(n349), .Z(n346) );
  GTECH_AND2 U386 ( .A(n168), .B(update_period[2]), .Z(n348) );
  GTECH_AND3 U387 ( .A(n350), .B(n351), .C(n349), .Z(n345) );
  GTECH_NAND2 U388 ( .A(n347), .B(n312), .Z(n349) );
  GTECH_NOT U389 ( .A(n167), .Z(n312) );
  GTECH_NOT U390 ( .A(update_period[3]), .Z(n347) );
  GTECH_OAI21 U391 ( .A(n352), .B(n320), .C(n175), .Z(n351) );
  GTECH_NOT U392 ( .A(n169), .Z(n320) );
  GTECH_OA21 U393 ( .A(n168), .B(update_period[2]), .C(n353), .Z(n350) );
  GTECH_OR_NOT U394 ( .A(n169), .B(n352), .Z(n353) );
  GTECH_NAND2 U395 ( .A(update_period[0]), .B(n170), .Z(n352) );
  GTECH_OA22 U396 ( .A(n162), .B(update_period[8]), .C(n161), .D(
        update_period[9]), .Z(n322) );
  GTECH_AO21 U397 ( .A(period[2]), .B(n214), .C(reset), .Z(N11) );
  GTECH_AO21 U398 ( .A(period[1]), .B(n214), .C(reset), .Z(N10) );
  GTECH_NOT U399 ( .A(n215), .Z(n214) );
  GTECH_NAND2 U400 ( .A(period_load), .B(n187), .Z(n215) );
  GTECH_NOT U401 ( .A(reset), .Z(n187) );
endmodule

