
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389;

  GTECH_MUX2 U142 ( .A(n281), .B(n282), .S(n283), .Z(sum[9]) );
  GTECH_XOR2 U143 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_XOR2 U144 ( .A(n284), .B(n286), .Z(n281) );
  GTECH_AO21 U145 ( .A(a[9]), .B(b[9]), .C(n287), .Z(n284) );
  GTECH_AO21 U146 ( .A(n288), .B(n283), .C(n289), .Z(sum[8]) );
  GTECH_MUX2 U147 ( .A(n290), .B(n291), .S(n292), .Z(sum[7]) );
  GTECH_NOT U148 ( .A(n293), .Z(n291) );
  GTECH_XOR2 U149 ( .A(n294), .B(n295), .Z(n293) );
  GTECH_AND2 U150 ( .A(n296), .B(n297), .Z(n295) );
  GTECH_AO21 U151 ( .A(n298), .B(n299), .C(n300), .Z(n297) );
  GTECH_XOR2 U152 ( .A(n294), .B(n301), .Z(n290) );
  GTECH_XOR2 U153 ( .A(a[7]), .B(b[7]), .Z(n294) );
  GTECH_OAI21 U154 ( .A(n302), .B(n296), .C(n303), .Z(sum[6]) );
  GTECH_MUX2 U155 ( .A(n304), .B(n305), .S(b[6]), .Z(n303) );
  GTECH_OR_NOT U156 ( .A(a[6]), .B(n302), .Z(n305) );
  GTECH_XOR2 U157 ( .A(n302), .B(a[6]), .Z(n304) );
  GTECH_AO21 U158 ( .A(n306), .B(n298), .C(n307), .Z(n302) );
  GTECH_NOT U159 ( .A(n308), .Z(n298) );
  GTECH_XOR2 U160 ( .A(n306), .B(n309), .Z(sum[5]) );
  GTECH_OR_NOT U161 ( .A(n308), .B(n310), .Z(n309) );
  GTECH_OAI2N2 U162 ( .A(b[4]), .B(a[4]), .C(n299), .D(n292), .Z(n306) );
  GTECH_NAND2 U163 ( .A(b[4]), .B(a[4]), .Z(n299) );
  GTECH_XOR2 U164 ( .A(n311), .B(n312), .Z(sum[4]) );
  GTECH_NOT U165 ( .A(n292), .Z(n311) );
  GTECH_MUX2 U166 ( .A(n313), .B(n314), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U167 ( .A(n315), .B(n316), .Z(n314) );
  GTECH_NOT U168 ( .A(n317), .Z(n313) );
  GTECH_XOR2 U169 ( .A(n315), .B(n318), .Z(n317) );
  GTECH_AND2 U170 ( .A(n319), .B(n320), .Z(n318) );
  GTECH_OAI21 U171 ( .A(b[2]), .B(a[2]), .C(n321), .Z(n319) );
  GTECH_XOR2 U172 ( .A(a[3]), .B(b[3]), .Z(n315) );
  GTECH_MUX2 U173 ( .A(n322), .B(n323), .S(n324), .Z(sum[2]) );
  GTECH_MUX2 U174 ( .A(n325), .B(n326), .S(n321), .Z(n323) );
  GTECH_AOI2N2 U175 ( .A(n327), .B(n328), .C(b[1]), .D(a[1]), .Z(n321) );
  GTECH_MUX2 U176 ( .A(n325), .B(n326), .S(n329), .Z(n322) );
  GTECH_OAI21 U177 ( .A(b[2]), .B(a[2]), .C(n320), .Z(n326) );
  GTECH_XOR2 U178 ( .A(a[2]), .B(b[2]), .Z(n325) );
  GTECH_MUX2 U179 ( .A(n330), .B(n331), .S(n332), .Z(sum[1]) );
  GTECH_XOR2 U180 ( .A(b[1]), .B(a[1]), .Z(n332) );
  GTECH_AO21 U181 ( .A(n324), .B(n328), .C(n333), .Z(n331) );
  GTECH_OAI21 U182 ( .A(n333), .B(n324), .C(n328), .Z(n330) );
  GTECH_NAND2 U183 ( .A(a[0]), .B(b[0]), .Z(n328) );
  GTECH_NOT U184 ( .A(cin), .Z(n324) );
  GTECH_MUX2 U185 ( .A(n334), .B(n335), .S(n336), .Z(sum[15]) );
  GTECH_XOR2 U186 ( .A(n337), .B(n338), .Z(n335) );
  GTECH_AND2 U187 ( .A(n339), .B(n340), .Z(n338) );
  GTECH_AO21 U188 ( .A(n341), .B(n342), .C(n343), .Z(n339) );
  GTECH_XOR2 U189 ( .A(n337), .B(n344), .Z(n334) );
  GTECH_XOR2 U190 ( .A(n345), .B(b[15]), .Z(n337) );
  GTECH_OAI21 U191 ( .A(n346), .B(n340), .C(n347), .Z(sum[14]) );
  GTECH_MUX2 U192 ( .A(n348), .B(n349), .S(b[14]), .Z(n347) );
  GTECH_OR_NOT U193 ( .A(a[14]), .B(n346), .Z(n349) );
  GTECH_XOR2 U194 ( .A(a[14]), .B(n346), .Z(n348) );
  GTECH_OA21 U195 ( .A(n350), .B(n336), .C(n343), .Z(n346) );
  GTECH_OA21 U196 ( .A(n351), .B(n352), .C(n353), .Z(n343) );
  GTECH_MUX2 U197 ( .A(n354), .B(n355), .S(n356), .Z(sum[13]) );
  GTECH_OA21 U198 ( .A(n336), .B(n357), .C(n352), .Z(n356) );
  GTECH_XOR2 U199 ( .A(b[13]), .B(a[13]), .Z(n355) );
  GTECH_OR_NOT U200 ( .A(n351), .B(n353), .Z(n354) );
  GTECH_AO21 U201 ( .A(n358), .B(n359), .C(n360), .Z(sum[12]) );
  GTECH_MUX2 U202 ( .A(n361), .B(n362), .S(n283), .Z(sum[11]) );
  GTECH_XOR2 U203 ( .A(n363), .B(n364), .Z(n362) );
  GTECH_NOT U204 ( .A(n365), .Z(n361) );
  GTECH_XOR2 U205 ( .A(n363), .B(n366), .Z(n365) );
  GTECH_AND2 U206 ( .A(n367), .B(n368), .Z(n366) );
  GTECH_OAI21 U207 ( .A(b[10]), .B(a[10]), .C(n369), .Z(n367) );
  GTECH_XOR2 U208 ( .A(a[11]), .B(b[11]), .Z(n363) );
  GTECH_OAI21 U209 ( .A(n370), .B(n368), .C(n371), .Z(sum[10]) );
  GTECH_MUX2 U210 ( .A(n372), .B(n373), .S(b[10]), .Z(n371) );
  GTECH_OR_NOT U211 ( .A(a[10]), .B(n370), .Z(n373) );
  GTECH_XOR2 U212 ( .A(a[10]), .B(n370), .Z(n372) );
  GTECH_AOI21 U213 ( .A(n374), .B(n283), .C(n369), .Z(n370) );
  GTECH_OAI2N2 U214 ( .A(n287), .B(n286), .C(a[9]), .D(b[9]), .Z(n369) );
  GTECH_XOR2 U215 ( .A(cin), .B(n375), .Z(sum[0]) );
  GTECH_AO21 U216 ( .A(n358), .B(n376), .C(n360), .Z(cout) );
  GTECH_AND_NOT U217 ( .A(n336), .B(n359), .Z(n360) );
  GTECH_OR_NOT U218 ( .A(n357), .B(n352), .Z(n359) );
  GTECH_NAND2 U219 ( .A(a[12]), .B(b[12]), .Z(n352) );
  GTECH_NOT U220 ( .A(n358), .Z(n336) );
  GTECH_OAI21 U221 ( .A(n344), .B(n345), .C(n377), .Z(n376) );
  GTECH_AO21 U222 ( .A(n345), .B(n344), .C(n378), .Z(n377) );
  GTECH_NOT U223 ( .A(b[15]), .Z(n378) );
  GTECH_NOT U224 ( .A(a[15]), .Z(n345) );
  GTECH_AND2 U225 ( .A(n379), .B(n340), .Z(n344) );
  GTECH_OR_NOT U226 ( .A(n341), .B(a[14]), .Z(n340) );
  GTECH_AO21 U227 ( .A(n342), .B(n341), .C(n350), .Z(n379) );
  GTECH_OA21 U228 ( .A(n357), .B(n351), .C(n353), .Z(n350) );
  GTECH_NAND2 U229 ( .A(b[13]), .B(a[13]), .Z(n353) );
  GTECH_NOR2 U230 ( .A(b[13]), .B(a[13]), .Z(n351) );
  GTECH_NOR2 U231 ( .A(b[12]), .B(a[12]), .Z(n357) );
  GTECH_NOT U232 ( .A(b[14]), .Z(n341) );
  GTECH_NOT U233 ( .A(a[14]), .Z(n342) );
  GTECH_AO21 U234 ( .A(n283), .B(n380), .C(n289), .Z(n358) );
  GTECH_NOR2 U235 ( .A(n283), .B(n288), .Z(n289) );
  GTECH_OR_NOT U236 ( .A(n285), .B(n286), .Z(n288) );
  GTECH_NAND2 U237 ( .A(b[8]), .B(a[8]), .Z(n286) );
  GTECH_OA21 U238 ( .A(a[11]), .B(n364), .C(n381), .Z(n380) );
  GTECH_AO21 U239 ( .A(n364), .B(a[11]), .C(b[11]), .Z(n381) );
  GTECH_NAND2 U240 ( .A(n382), .B(n368), .Z(n364) );
  GTECH_NAND2 U241 ( .A(b[10]), .B(a[10]), .Z(n368) );
  GTECH_OAI21 U242 ( .A(a[10]), .B(b[10]), .C(n374), .Z(n382) );
  GTECH_OAI2N2 U243 ( .A(n285), .B(n287), .C(a[9]), .D(b[9]), .Z(n374) );
  GTECH_NOR2 U244 ( .A(b[9]), .B(a[9]), .Z(n287) );
  GTECH_NOR2 U245 ( .A(a[8]), .B(b[8]), .Z(n285) );
  GTECH_MUX2 U246 ( .A(n383), .B(n312), .S(n292), .Z(n283) );
  GTECH_MUX2 U247 ( .A(n384), .B(n385), .S(cin), .Z(n292) );
  GTECH_AOI21 U248 ( .A(n316), .B(a[3]), .C(n386), .Z(n385) );
  GTECH_OA21 U249 ( .A(a[3]), .B(n316), .C(b[3]), .Z(n386) );
  GTECH_NAND2 U250 ( .A(n320), .B(n387), .Z(n316) );
  GTECH_OAI21 U251 ( .A(a[2]), .B(b[2]), .C(n329), .Z(n387) );
  GTECH_AOI2N2 U252 ( .A(n327), .B(n333), .C(b[1]), .D(a[1]), .Z(n329) );
  GTECH_NOR2 U253 ( .A(a[0]), .B(b[0]), .Z(n333) );
  GTECH_NAND2 U254 ( .A(a[1]), .B(b[1]), .Z(n327) );
  GTECH_NAND2 U255 ( .A(b[2]), .B(a[2]), .Z(n320) );
  GTECH_NOT U256 ( .A(n375), .Z(n384) );
  GTECH_XOR2 U257 ( .A(a[0]), .B(b[0]), .Z(n375) );
  GTECH_XOR2 U258 ( .A(a[4]), .B(b[4]), .Z(n312) );
  GTECH_OA21 U259 ( .A(a[7]), .B(n301), .C(n388), .Z(n383) );
  GTECH_AO21 U260 ( .A(n301), .B(a[7]), .C(b[7]), .Z(n388) );
  GTECH_OAI21 U261 ( .A(n389), .B(n300), .C(n296), .Z(n301) );
  GTECH_NAND2 U262 ( .A(b[6]), .B(a[6]), .Z(n296) );
  GTECH_OAI21 U263 ( .A(b[6]), .B(a[6]), .C(n310), .Z(n300) );
  GTECH_NOT U264 ( .A(n307), .Z(n310) );
  GTECH_NOR2 U265 ( .A(b[5]), .B(a[5]), .Z(n307) );
  GTECH_NOR3 U266 ( .A(a[4]), .B(b[4]), .C(n308), .Z(n389) );
  GTECH_AND2 U267 ( .A(a[5]), .B(b[5]), .Z(n308) );
endmodule

