
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364;

  GTECH_MUX2 U128 ( .A(n267), .B(n268), .S(n269), .Z(sum[9]) );
  GTECH_XOR2 U129 ( .A(n270), .B(n271), .Z(n268) );
  GTECH_XOR2 U130 ( .A(n271), .B(n272), .Z(n267) );
  GTECH_AO21 U131 ( .A(a[9]), .B(b[9]), .C(n273), .Z(n271) );
  GTECH_XNOR2 U132 ( .A(n274), .B(n269), .Z(sum[8]) );
  GTECH_MUX2 U133 ( .A(n275), .B(n276), .S(n277), .Z(sum[7]) );
  GTECH_XOR2 U134 ( .A(n278), .B(n279), .Z(n276) );
  GTECH_XNOR2 U135 ( .A(n278), .B(n280), .Z(n275) );
  GTECH_AOI22 U136 ( .A(n281), .B(n282), .C(a[6]), .D(b[6]), .Z(n280) );
  GTECH_XOR2 U137 ( .A(a[7]), .B(b[7]), .Z(n278) );
  GTECH_MUX2 U138 ( .A(n283), .B(n284), .S(n277), .Z(sum[6]) );
  GTECH_XNOR2 U139 ( .A(n285), .B(n286), .Z(n284) );
  GTECH_XNOR2 U140 ( .A(n281), .B(n286), .Z(n283) );
  GTECH_AO21 U141 ( .A(a[6]), .B(b[6]), .C(n287), .Z(n286) );
  GTECH_NOT U142 ( .A(n282), .Z(n287) );
  GTECH_AO21 U143 ( .A(n288), .B(n289), .C(n290), .Z(n281) );
  GTECH_MUX2 U144 ( .A(n291), .B(n292), .S(n293), .Z(sum[5]) );
  GTECH_AND_NOT U145 ( .A(n288), .B(n290), .Z(n293) );
  GTECH_OAI21 U146 ( .A(n289), .B(n277), .C(n294), .Z(n292) );
  GTECH_AO21 U147 ( .A(n294), .B(n277), .C(n289), .Z(n291) );
  GTECH_XOR2 U148 ( .A(n277), .B(n295), .Z(sum[4]) );
  GTECH_MUX2 U149 ( .A(n296), .B(n297), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U150 ( .A(n298), .B(n299), .Z(n297) );
  GTECH_XNOR2 U151 ( .A(n298), .B(n300), .Z(n296) );
  GTECH_AOI22 U152 ( .A(n301), .B(n302), .C(a[2]), .D(b[2]), .Z(n300) );
  GTECH_XOR2 U153 ( .A(a[3]), .B(b[3]), .Z(n298) );
  GTECH_MUX2 U154 ( .A(n303), .B(n304), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U155 ( .A(n305), .B(n306), .Z(n304) );
  GTECH_XNOR2 U156 ( .A(n302), .B(n306), .Z(n303) );
  GTECH_AO21 U157 ( .A(a[2]), .B(b[2]), .C(n307), .Z(n306) );
  GTECH_NOT U158 ( .A(n301), .Z(n307) );
  GTECH_AO21 U159 ( .A(n308), .B(n309), .C(n310), .Z(n302) );
  GTECH_AO22 U160 ( .A(n311), .B(n312), .C(n313), .D(n314), .Z(sum[1]) );
  GTECH_OAI21 U161 ( .A(cin), .B(n309), .C(n315), .Z(n314) );
  GTECH_XOR2 U162 ( .A(b[1]), .B(a[1]), .Z(n313) );
  GTECH_OAI21 U163 ( .A(n316), .B(n317), .C(n318), .Z(n312) );
  GTECH_NOT U164 ( .A(n309), .Z(n318) );
  GTECH_OR_NOT U165 ( .A(n310), .B(n308), .Z(n311) );
  GTECH_MUX2 U166 ( .A(n319), .B(n320), .S(n321), .Z(sum[15]) );
  GTECH_XNOR2 U167 ( .A(n322), .B(n323), .Z(n320) );
  GTECH_AOI22 U168 ( .A(a[14]), .B(b[14]), .C(n324), .D(n325), .Z(n323) );
  GTECH_XOR2 U169 ( .A(n322), .B(n326), .Z(n319) );
  GTECH_XOR2 U170 ( .A(a[15]), .B(b[15]), .Z(n322) );
  GTECH_MUX2 U171 ( .A(n327), .B(n328), .S(n321), .Z(sum[14]) );
  GTECH_XNOR2 U172 ( .A(n325), .B(n329), .Z(n328) );
  GTECH_OAI2N2 U173 ( .A(n330), .B(n331), .C(a[13]), .D(b[13]), .Z(n325) );
  GTECH_XNOR2 U174 ( .A(n332), .B(n329), .Z(n327) );
  GTECH_AO21 U175 ( .A(a[14]), .B(b[14]), .C(n333), .Z(n329) );
  GTECH_NOT U176 ( .A(n324), .Z(n333) );
  GTECH_MUX2 U177 ( .A(n334), .B(n335), .S(n321), .Z(sum[13]) );
  GTECH_XOR2 U178 ( .A(n336), .B(n331), .Z(n335) );
  GTECH_XNOR2 U179 ( .A(n337), .B(n336), .Z(n334) );
  GTECH_AO21 U180 ( .A(a[13]), .B(b[13]), .C(n330), .Z(n336) );
  GTECH_NAND2 U181 ( .A(n338), .B(n339), .Z(sum[12]) );
  GTECH_AO21 U182 ( .A(n331), .B(n337), .C(n321), .Z(n339) );
  GTECH_MUX2 U183 ( .A(n340), .B(n341), .S(n269), .Z(sum[11]) );
  GTECH_XOR2 U184 ( .A(n342), .B(n343), .Z(n341) );
  GTECH_XNOR2 U185 ( .A(n342), .B(n344), .Z(n340) );
  GTECH_AOI22 U186 ( .A(a[10]), .B(b[10]), .C(n345), .D(n346), .Z(n344) );
  GTECH_XOR2 U187 ( .A(a[11]), .B(b[11]), .Z(n342) );
  GTECH_MUX2 U188 ( .A(n347), .B(n348), .S(n269), .Z(sum[10]) );
  GTECH_XNOR2 U189 ( .A(n349), .B(n350), .Z(n348) );
  GTECH_XNOR2 U190 ( .A(n346), .B(n350), .Z(n347) );
  GTECH_AO21 U191 ( .A(a[10]), .B(b[10]), .C(n351), .Z(n350) );
  GTECH_NOT U192 ( .A(n345), .Z(n351) );
  GTECH_OAI2N2 U193 ( .A(n273), .B(n272), .C(a[9]), .D(b[9]), .Z(n346) );
  GTECH_NOT U194 ( .A(n352), .Z(n272) );
  GTECH_NAND2 U195 ( .A(n353), .B(n354), .Z(sum[0]) );
  GTECH_OAI21 U196 ( .A(n309), .B(n316), .C(cin), .Z(n354) );
  GTECH_OAI21 U197 ( .A(n355), .B(n321), .C(n338), .Z(cout) );
  GTECH_NAND3 U198 ( .A(n331), .B(n337), .C(n321), .Z(n338) );
  GTECH_NAND2 U199 ( .A(b[12]), .B(a[12]), .Z(n331) );
  GTECH_MUX2 U200 ( .A(n274), .B(n356), .S(n269), .Z(n321) );
  GTECH_MUX2 U201 ( .A(n295), .B(n357), .S(n277), .Z(n269) );
  GTECH_OAI21 U202 ( .A(n358), .B(n317), .C(n353), .Z(n277) );
  GTECH_OR3 U203 ( .A(n309), .B(cin), .C(n316), .Z(n353) );
  GTECH_AND2 U204 ( .A(b[0]), .B(a[0]), .Z(n309) );
  GTECH_NOT U205 ( .A(cin), .Z(n317) );
  GTECH_AOI2N2 U206 ( .A(n359), .B(b[3]), .C(n299), .D(n360), .Z(n358) );
  GTECH_NOT U207 ( .A(a[3]), .Z(n360) );
  GTECH_OR_NOT U208 ( .A(a[3]), .B(n299), .Z(n359) );
  GTECH_AOI22 U209 ( .A(n305), .B(n301), .C(a[2]), .D(b[2]), .Z(n299) );
  GTECH_OR2 U210 ( .A(a[2]), .B(b[2]), .Z(n301) );
  GTECH_AO21 U211 ( .A(n315), .B(n308), .C(n310), .Z(n305) );
  GTECH_AND2 U212 ( .A(b[1]), .B(a[1]), .Z(n310) );
  GTECH_OR2 U213 ( .A(b[1]), .B(a[1]), .Z(n308) );
  GTECH_NOT U214 ( .A(n316), .Z(n315) );
  GTECH_NOR2 U215 ( .A(a[0]), .B(b[0]), .Z(n316) );
  GTECH_AO22 U216 ( .A(n279), .B(a[7]), .C(n361), .D(b[7]), .Z(n357) );
  GTECH_OR2 U217 ( .A(a[7]), .B(n279), .Z(n361) );
  GTECH_AO22 U218 ( .A(n285), .B(n282), .C(a[6]), .D(b[6]), .Z(n279) );
  GTECH_OR2 U219 ( .A(a[6]), .B(b[6]), .Z(n282) );
  GTECH_AO21 U220 ( .A(n294), .B(n288), .C(n290), .Z(n285) );
  GTECH_AND2 U221 ( .A(b[5]), .B(a[5]), .Z(n290) );
  GTECH_OR2 U222 ( .A(a[5]), .B(b[5]), .Z(n288) );
  GTECH_AND_NOT U223 ( .A(n294), .B(n289), .Z(n295) );
  GTECH_AND2 U224 ( .A(b[4]), .B(a[4]), .Z(n289) );
  GTECH_OR2 U225 ( .A(a[4]), .B(b[4]), .Z(n294) );
  GTECH_AOI22 U226 ( .A(n343), .B(a[11]), .C(n362), .D(b[11]), .Z(n356) );
  GTECH_OR2 U227 ( .A(a[11]), .B(n343), .Z(n362) );
  GTECH_AO22 U228 ( .A(a[10]), .B(b[10]), .C(n349), .D(n345), .Z(n343) );
  GTECH_OR2 U229 ( .A(a[10]), .B(b[10]), .Z(n345) );
  GTECH_OAI2N2 U230 ( .A(n270), .B(n273), .C(a[9]), .D(b[9]), .Z(n349) );
  GTECH_NOR2 U231 ( .A(a[9]), .B(b[9]), .Z(n273) );
  GTECH_OR2 U232 ( .A(n270), .B(n352), .Z(n274) );
  GTECH_AND2 U233 ( .A(b[8]), .B(a[8]), .Z(n352) );
  GTECH_NOR2 U234 ( .A(a[8]), .B(b[8]), .Z(n270) );
  GTECH_AOI22 U235 ( .A(n326), .B(a[15]), .C(n363), .D(b[15]), .Z(n355) );
  GTECH_OR2 U236 ( .A(n326), .B(a[15]), .Z(n363) );
  GTECH_AO22 U237 ( .A(a[14]), .B(b[14]), .C(n332), .D(n324), .Z(n326) );
  GTECH_OR2 U238 ( .A(a[14]), .B(b[14]), .Z(n324) );
  GTECH_AO22 U239 ( .A(n337), .B(n364), .C(a[13]), .D(b[13]), .Z(n332) );
  GTECH_NOT U240 ( .A(n330), .Z(n364) );
  GTECH_NOR2 U241 ( .A(a[13]), .B(b[13]), .Z(n330) );
  GTECH_OR2 U242 ( .A(a[12]), .B(b[12]), .Z(n337) );
endmodule

