
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394;

  GTECH_MUX2 U144 ( .A(n283), .B(n284), .S(n285), .Z(sum[9]) );
  GTECH_XNOR2 U145 ( .A(n286), .B(n287), .Z(n284) );
  GTECH_XNOR2 U146 ( .A(n288), .B(n287), .Z(n283) );
  GTECH_AOI21 U147 ( .A(a[9]), .B(b[9]), .C(n289), .Z(n287) );
  GTECH_NAND2 U148 ( .A(n290), .B(n291), .Z(sum[8]) );
  GTECH_AO21 U149 ( .A(n288), .B(n292), .C(n293), .Z(n290) );
  GTECH_MUX2 U150 ( .A(n294), .B(n295), .S(n296), .Z(sum[7]) );
  GTECH_XNOR2 U151 ( .A(n297), .B(n298), .Z(n295) );
  GTECH_AND2 U152 ( .A(n299), .B(n300), .Z(n297) );
  GTECH_AO21 U153 ( .A(n301), .B(n302), .C(n303), .Z(n300) );
  GTECH_ADD_AB U154 ( .A(n304), .B(n298), .S(n294) );
  GTECH_ADD_AB U155 ( .A(b[7]), .B(a[7]), .S(n298) );
  GTECH_OAI21 U156 ( .A(n305), .B(n299), .C(n306), .Z(sum[6]) );
  GTECH_MUX2 U157 ( .A(n307), .B(n308), .S(b[6]), .Z(n306) );
  GTECH_NAND2 U158 ( .A(n302), .B(n305), .Z(n308) );
  GTECH_XNOR2 U159 ( .A(n302), .B(n305), .Z(n307) );
  GTECH_OA21 U160 ( .A(n309), .B(n296), .C(n303), .Z(n305) );
  GTECH_OAI21 U161 ( .A(n310), .B(n311), .C(n312), .Z(n303) );
  GTECH_MUX2 U162 ( .A(n313), .B(n314), .S(n315), .Z(sum[5]) );
  GTECH_AND_NOT U163 ( .A(n312), .B(n310), .Z(n315) );
  GTECH_OAI21 U164 ( .A(a[4]), .B(n316), .C(n317), .Z(n314) );
  GTECH_AO21 U165 ( .A(n316), .B(a[4]), .C(b[4]), .Z(n317) );
  GTECH_AO21 U166 ( .A(n318), .B(n316), .C(n311), .Z(n313) );
  GTECH_ADD_AB U167 ( .A(n319), .B(n296), .S(sum[4]) );
  GTECH_MUX2 U168 ( .A(n320), .B(n321), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U169 ( .A(n322), .B(n323), .Z(n321) );
  GTECH_ADD_AB U170 ( .A(n324), .B(n323), .S(n320) );
  GTECH_XNOR2 U171 ( .A(b[3]), .B(a[3]), .Z(n323) );
  GTECH_AND2 U172 ( .A(n325), .B(n326), .Z(n324) );
  GTECH_AO21 U173 ( .A(n327), .B(n328), .C(n329), .Z(n326) );
  GTECH_MUX2 U174 ( .A(n330), .B(n331), .S(n332), .Z(sum[2]) );
  GTECH_MUX2 U175 ( .A(n333), .B(n334), .S(n329), .Z(n331) );
  GTECH_AO21 U176 ( .A(n335), .B(n336), .C(n337), .Z(n329) );
  GTECH_MUX2 U177 ( .A(n334), .B(n333), .S(n338), .Z(n330) );
  GTECH_OAI21 U178 ( .A(b[2]), .B(a[2]), .C(n325), .Z(n333) );
  GTECH_ADD_AB U179 ( .A(n327), .B(n328), .S(n334) );
  GTECH_NOT U180 ( .A(a[2]), .Z(n328) );
  GTECH_MUX2 U181 ( .A(n339), .B(n340), .S(n341), .Z(sum[1]) );
  GTECH_AND_NOT U182 ( .A(n335), .B(n337), .Z(n341) );
  GTECH_AO21 U183 ( .A(n332), .B(n336), .C(n342), .Z(n340) );
  GTECH_OAI21 U184 ( .A(n342), .B(n332), .C(n336), .Z(n339) );
  GTECH_NAND2 U185 ( .A(b[0]), .B(a[0]), .Z(n336) );
  GTECH_NOT U186 ( .A(cin), .Z(n332) );
  GTECH_MUX2 U187 ( .A(n343), .B(n344), .S(n345), .Z(sum[15]) );
  GTECH_XNOR2 U188 ( .A(n346), .B(n347), .Z(n344) );
  GTECH_OA21 U189 ( .A(n348), .B(n349), .C(n350), .Z(n346) );
  GTECH_ADD_AB U190 ( .A(n351), .B(n347), .S(n343) );
  GTECH_ADD_AB U191 ( .A(b[15]), .B(a[15]), .S(n347) );
  GTECH_MUX2 U192 ( .A(n352), .B(n353), .S(n354), .Z(sum[14]) );
  GTECH_OA21 U193 ( .A(n355), .B(n345), .C(n349), .Z(n354) );
  GTECH_AND2 U194 ( .A(n356), .B(n357), .Z(n349) );
  GTECH_OAI21 U195 ( .A(b[13]), .B(a[13]), .C(n358), .Z(n356) );
  GTECH_ADD_AB U196 ( .A(b[14]), .B(a[14]), .S(n353) );
  GTECH_OR_NOT U197 ( .A(n348), .B(n350), .Z(n352) );
  GTECH_MUX2 U198 ( .A(n359), .B(n360), .S(n345), .Z(sum[13]) );
  GTECH_ADD_AB U199 ( .A(n358), .B(n361), .S(n360) );
  GTECH_ADD_AB U200 ( .A(n362), .B(n361), .S(n359) );
  GTECH_OA21 U201 ( .A(a[13]), .B(b[13]), .C(n357), .Z(n361) );
  GTECH_NAND2 U202 ( .A(n363), .B(n364), .Z(sum[12]) );
  GTECH_OAI21 U203 ( .A(n358), .B(n365), .C(n366), .Z(n363) );
  GTECH_MUX2 U204 ( .A(n367), .B(n368), .S(n285), .Z(sum[11]) );
  GTECH_ADD_AB U205 ( .A(n369), .B(n370), .S(n368) );
  GTECH_XNOR2 U206 ( .A(n371), .B(n370), .Z(n367) );
  GTECH_ADD_AB U207 ( .A(b[11]), .B(a[11]), .S(n370) );
  GTECH_AND2 U208 ( .A(n372), .B(n373), .Z(n371) );
  GTECH_OAI21 U209 ( .A(b[10]), .B(a[10]), .C(n374), .Z(n373) );
  GTECH_OAI21 U210 ( .A(n375), .B(n372), .C(n376), .Z(sum[10]) );
  GTECH_MUX2 U211 ( .A(n377), .B(n378), .S(b[10]), .Z(n376) );
  GTECH_OR_NOT U212 ( .A(a[10]), .B(n375), .Z(n378) );
  GTECH_ADD_AB U213 ( .A(a[10]), .B(n375), .S(n377) );
  GTECH_AOI21 U214 ( .A(n379), .B(n285), .C(n374), .Z(n375) );
  GTECH_OAI2N2 U215 ( .A(n289), .B(n288), .C(a[9]), .D(b[9]), .Z(n374) );
  GTECH_NOT U216 ( .A(n293), .Z(n285) );
  GTECH_ADD_AB U217 ( .A(cin), .B(n380), .S(sum[0]) );
  GTECH_OAI21 U218 ( .A(n345), .B(n381), .C(n364), .Z(cout) );
  GTECH_OR3 U219 ( .A(n358), .B(n365), .C(n366), .Z(n364) );
  GTECH_AND2 U220 ( .A(a[12]), .B(b[12]), .Z(n358) );
  GTECH_AOI21 U221 ( .A(n351), .B(a[15]), .C(n382), .Z(n381) );
  GTECH_OA21 U222 ( .A(a[15]), .B(n351), .C(b[15]), .Z(n382) );
  GTECH_NAND2 U223 ( .A(n383), .B(n350), .Z(n351) );
  GTECH_NAND2 U224 ( .A(a[14]), .B(b[14]), .Z(n350) );
  GTECH_AO21 U225 ( .A(n355), .B(n357), .C(n348), .Z(n383) );
  GTECH_NOR2 U226 ( .A(a[14]), .B(b[14]), .Z(n348) );
  GTECH_NAND2 U227 ( .A(b[13]), .B(a[13]), .Z(n357) );
  GTECH_OAI21 U228 ( .A(b[13]), .B(a[13]), .C(n362), .Z(n355) );
  GTECH_NOT U229 ( .A(n365), .Z(n362) );
  GTECH_NOR2 U230 ( .A(b[12]), .B(a[12]), .Z(n365) );
  GTECH_NOT U231 ( .A(n366), .Z(n345) );
  GTECH_OAI21 U232 ( .A(n384), .B(n293), .C(n291), .Z(n366) );
  GTECH_NAND3 U233 ( .A(n288), .B(n292), .C(n293), .Z(n291) );
  GTECH_NOT U234 ( .A(n286), .Z(n292) );
  GTECH_NAND2 U235 ( .A(b[8]), .B(a[8]), .Z(n288) );
  GTECH_MUX2 U236 ( .A(n385), .B(n319), .S(n296), .Z(n293) );
  GTECH_NOT U237 ( .A(n316), .Z(n296) );
  GTECH_MUX2 U238 ( .A(n380), .B(n386), .S(cin), .Z(n316) );
  GTECH_OA21 U239 ( .A(a[3]), .B(n322), .C(n387), .Z(n386) );
  GTECH_AO21 U240 ( .A(n322), .B(a[3]), .C(b[3]), .Z(n387) );
  GTECH_NAND2 U241 ( .A(n388), .B(n325), .Z(n322) );
  GTECH_OR_NOT U242 ( .A(n327), .B(a[2]), .Z(n325) );
  GTECH_NOT U243 ( .A(b[2]), .Z(n327) );
  GTECH_OAI21 U244 ( .A(a[2]), .B(b[2]), .C(n338), .Z(n388) );
  GTECH_AOI21 U245 ( .A(n335), .B(n342), .C(n337), .Z(n338) );
  GTECH_NOR2 U246 ( .A(b[1]), .B(a[1]), .Z(n337) );
  GTECH_AND_NOT U247 ( .A(n389), .B(b[0]), .Z(n342) );
  GTECH_NAND2 U248 ( .A(b[1]), .B(a[1]), .Z(n335) );
  GTECH_ADD_AB U249 ( .A(n390), .B(n389), .S(n380) );
  GTECH_NOT U250 ( .A(a[0]), .Z(n389) );
  GTECH_NOT U251 ( .A(b[0]), .Z(n390) );
  GTECH_OR_NOT U252 ( .A(n311), .B(n318), .Z(n319) );
  GTECH_AND2 U253 ( .A(a[4]), .B(b[4]), .Z(n311) );
  GTECH_AOI21 U254 ( .A(n304), .B(a[7]), .C(n391), .Z(n385) );
  GTECH_OA21 U255 ( .A(a[7]), .B(n304), .C(b[7]), .Z(n391) );
  GTECH_NAND2 U256 ( .A(n392), .B(n299), .Z(n304) );
  GTECH_OR_NOT U257 ( .A(n302), .B(b[6]), .Z(n299) );
  GTECH_AO21 U258 ( .A(n302), .B(n301), .C(n309), .Z(n392) );
  GTECH_OAI21 U259 ( .A(n310), .B(n318), .C(n312), .Z(n309) );
  GTECH_OR2 U260 ( .A(a[5]), .B(b[5]), .Z(n312) );
  GTECH_OR2 U261 ( .A(a[4]), .B(b[4]), .Z(n318) );
  GTECH_AND2 U262 ( .A(b[5]), .B(a[5]), .Z(n310) );
  GTECH_NOT U263 ( .A(b[6]), .Z(n301) );
  GTECH_NOT U264 ( .A(a[6]), .Z(n302) );
  GTECH_AOI21 U265 ( .A(n369), .B(a[11]), .C(n393), .Z(n384) );
  GTECH_OA21 U266 ( .A(a[11]), .B(n369), .C(b[11]), .Z(n393) );
  GTECH_NAND2 U267 ( .A(n394), .B(n372), .Z(n369) );
  GTECH_NAND2 U268 ( .A(a[10]), .B(b[10]), .Z(n372) );
  GTECH_OAI21 U269 ( .A(a[10]), .B(b[10]), .C(n379), .Z(n394) );
  GTECH_OAI2N2 U270 ( .A(n286), .B(n289), .C(a[9]), .D(b[9]), .Z(n379) );
  GTECH_NOR2 U271 ( .A(a[9]), .B(b[9]), .Z(n289) );
  GTECH_NOR2 U272 ( .A(a[8]), .B(b[8]), .Z(n286) );
endmodule

