
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(1'b0), .K(1'b0), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n249) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(1'b0), .K(1'b0), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(1'b0), .K(1'b0), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(1'b0), .K(1'b0), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(1'b0), .K(1'b0), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(1'b0), .K(1'b0), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]) );
  GTECH_FJK1S A_reg_15_ ( .J(1'b0), .K(1'b0), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n265) );
  GTECH_FJK1S A_reg_14_ ( .J(1'b0), .K(1'b0), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n264) );
  GTECH_FJK1S A_reg_13_ ( .J(1'b0), .K(1'b0), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n263) );
  GTECH_FJK1S A_reg_12_ ( .J(1'b0), .K(1'b0), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n262) );
  GTECH_FJK1S A_reg_11_ ( .J(1'b0), .K(1'b0), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n261) );
  GTECH_FJK1S A_reg_10_ ( .J(1'b0), .K(1'b0), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n260) );
  GTECH_FJK1S A_reg_9_ ( .J(1'b0), .K(1'b0), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n259) );
  GTECH_FJK1S A_reg_8_ ( .J(1'b0), .K(1'b0), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n258) );
  GTECH_FJK1S A_reg_7_ ( .J(1'b0), .K(1'b0), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n257) );
  GTECH_FJK1S A_reg_6_ ( .J(1'b0), .K(1'b0), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n256) );
  GTECH_FJK1S A_reg_5_ ( .J(1'b0), .K(1'b0), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n255) );
  GTECH_FJK1S A_reg_4_ ( .J(1'b0), .K(1'b0), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n254) );
  GTECH_FJK1S A_reg_3_ ( .J(1'b0), .K(1'b0), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n253) );
  GTECH_FJK1S A_reg_2_ ( .J(1'b0), .K(1'b0), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n252) );
  GTECH_FJK1S A_reg_1_ ( .J(1'b0), .K(1'b0), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n251) );
  GTECH_FJK1S A_reg_0_ ( .J(1'b0), .K(1'b0), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n250) );
  GTECH_FJK1S Prod_reg_0_ ( .J(1'b0), .K(1'b0), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(1'b0), .K(1'b0), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(1'b0), .K(1'b0), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(1'b0), .K(1'b0), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(1'b0), .K(1'b0), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(1'b0), .K(1'b0), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(1'b0), .K(1'b0), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(1'b0), .K(1'b0), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(1'b0), .K(1'b0), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(1'b0), .K(1'b0), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(1'b0), .K(1'b0), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(1'b0), .K(1'b0), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(1'b0), .K(1'b0), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(1'b0), .K(1'b0), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(1'b0), .K(1'b0), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(1'b0), .K(1'b0), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(1'b0), .K(1'b0), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(1'b0), .K(1'b0), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(1'b0), .K(1'b0), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(1'b0), .K(1'b0), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(1'b0), .K(1'b0), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(1'b0), .K(1'b0), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(1'b0), .K(1'b0), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(1'b0), .K(1'b0), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(1'b0), .K(1'b0), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(1'b0), .K(1'b0), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(1'b0), .K(1'b0), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(1'b0), .K(1'b0), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(1'b0), .K(1'b0), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(1'b0), .K(1'b0), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(1'b0), .K(1'b0), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(1'b0), .K(1'b0), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(1'b0), .K(1'b0), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(1'b0), .K(1'b0), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(1'b0), .K(1'b0), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(1'b0), .K(1'b0), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(1'b0), .K(1'b0), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(1'b0), .K(1'b0), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(1'b0), .K(1'b0), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(1'b0), .K(1'b0), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(1'b0), .K(1'b0), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(1'b0), .K(1'b0), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(1'b0), .K(1'b0), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(1'b0), .K(1'b0), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(1'b0), .K(1'b0), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(1'b0), .K(1'b0), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(1'b0), .K(1'b0), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(1'b0), .K(1'b0), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(1'b0), .K(1'b0), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(1'b0), .K(1'b0), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(1'b0), .K(1'b0), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(1'b0), .K(1'b0), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(1'b0), .K(1'b0), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(1'b0), .K(1'b0), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(1'b0), .K(1'b0), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(1'b0), .K(1'b0), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(1'b0), .K(1'b0), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(1'b0), .K(1'b0), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(1'b0), .K(1'b0), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(1'b0), .K(1'b0), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(1'b0), .K(1'b0), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(1'b0), .K(1'b0), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(1'b0), .K(1'b0), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(1'b0), .K(1'b0), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(1'b0), .K(1'b0), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(1'b0), .K(1'b0), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_NOT U251 ( .A(n267), .Z(N99) );
  GTECH_AOI222 U252 ( .A(n268), .B(n269), .C(n270), .D(n271), .E(n272), .F(
        n273), .Z(n267) );
  GTECH_NOT U253 ( .A(n274), .Z(N98) );
  GTECH_AOI222 U254 ( .A(n270), .B(n275), .C(n276), .D(n277), .E(R[15]), .F(
        n278), .Z(n274) );
  GTECH_NAND2 U255 ( .A(n279), .B(n280), .Z(n276) );
  GTECH_OAI2N2 U256 ( .A(n13), .B(n281), .C(R[14]), .D(n278), .Z(N97) );
  GTECH_OAI2N2 U257 ( .A(n14), .B(n281), .C(R[13]), .D(n278), .Z(N96) );
  GTECH_OAI2N2 U258 ( .A(n15), .B(n281), .C(R[12]), .D(n278), .Z(N95) );
  GTECH_OAI2N2 U259 ( .A(n16), .B(n281), .C(R[11]), .D(n278), .Z(N94) );
  GTECH_OAI2N2 U260 ( .A(n17), .B(n281), .C(R[10]), .D(n278), .Z(N93) );
  GTECH_OAI2N2 U261 ( .A(n18), .B(n281), .C(R[9]), .D(n278), .Z(N92) );
  GTECH_OAI2N2 U262 ( .A(n19), .B(n281), .C(R[8]), .D(n278), .Z(N91) );
  GTECH_OAI2N2 U263 ( .A(n20), .B(n281), .C(R[7]), .D(n278), .Z(N90) );
  GTECH_OAI2N2 U264 ( .A(n21), .B(n281), .C(R[6]), .D(n278), .Z(N89) );
  GTECH_OAI2N2 U265 ( .A(n22), .B(n281), .C(R[5]), .D(n278), .Z(N88) );
  GTECH_OAI2N2 U266 ( .A(n23), .B(n281), .C(R[4]), .D(n278), .Z(N87) );
  GTECH_OAI2N2 U267 ( .A(n24), .B(n281), .C(R[3]), .D(n278), .Z(N86) );
  GTECH_OAI2N2 U268 ( .A(n25), .B(n281), .C(R[2]), .D(n278), .Z(N85) );
  GTECH_OAI2N2 U269 ( .A(n26), .B(n281), .C(R[1]), .D(n278), .Z(N84) );
  GTECH_OAI2N2 U270 ( .A(n27), .B(n281), .C(R[0]), .D(n278), .Z(N83) );
  GTECH_AND2 U271 ( .A(M[15]), .B(n278), .Z(N42) );
  GTECH_AND2 U272 ( .A(M[14]), .B(n278), .Z(N39) );
  GTECH_AND2 U273 ( .A(M[13]), .B(n278), .Z(N38) );
  GTECH_AND2 U274 ( .A(M[12]), .B(n278), .Z(N37) );
  GTECH_AND2 U275 ( .A(M[11]), .B(n278), .Z(N36) );
  GTECH_AND2 U276 ( .A(M[10]), .B(n278), .Z(N35) );
  GTECH_AND2 U277 ( .A(M[9]), .B(n278), .Z(N34) );
  GTECH_AND2 U278 ( .A(M[8]), .B(n278), .Z(N33) );
  GTECH_AND2 U279 ( .A(M[7]), .B(n278), .Z(N32) );
  GTECH_AND2 U280 ( .A(M[6]), .B(n278), .Z(N31) );
  GTECH_AND2 U281 ( .A(M[5]), .B(n278), .Z(N30) );
  GTECH_AND2 U282 ( .A(M[4]), .B(n278), .Z(N29) );
  GTECH_AND2 U283 ( .A(M[3]), .B(n278), .Z(N28) );
  GTECH_AND2 U284 ( .A(M[2]), .B(n278), .Z(N27) );
  GTECH_AND2 U285 ( .A(M[1]), .B(n278), .Z(N26) );
  GTECH_AND2 U286 ( .A(M[0]), .B(n278), .Z(N25) );
  GTECH_NOT U287 ( .A(n282), .Z(n278) );
  GTECH_NAND2 U288 ( .A(n282), .B(n283), .Z(N19) );
  GTECH_NAND3 U289 ( .A(n284), .B(n285), .C(n286), .Z(n283) );
  GTECH_NAND3 U290 ( .A(n287), .B(n288), .C(n281), .Z(N18) );
  GTECH_AND2 U291 ( .A(n286), .B(n289), .Z(N17) );
  GTECH_OAI21 U292 ( .A(n8), .B(n290), .C(n284), .Z(n289) );
  GTECH_AND2 U293 ( .A(n286), .B(n291), .Z(N16) );
  GTECH_OAI21 U294 ( .A(n7), .B(n292), .C(n293), .Z(n291) );
  GTECH_NOT U295 ( .A(n294), .Z(N152) );
  GTECH_AOI222 U296 ( .A(n295), .B(n296), .C(n297), .D(n298), .E(n299), .F(
        n300), .Z(n294) );
  GTECH_NAND2 U297 ( .A(n288), .B(n301), .Z(N151) );
  GTECH_NOT U298 ( .A(n302), .Z(N150) );
  GTECH_AOI222 U299 ( .A(n303), .B(n295), .C(n297), .D(n304), .E(n299), .F(
        n305), .Z(n302) );
  GTECH_MUX2 U300 ( .A(n306), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND_NOT U301 ( .A(n286), .B(n249), .Z(n306) );
  GTECH_NOT U302 ( .A(n307), .Z(N149) );
  GTECH_AOI222 U303 ( .A(n308), .B(n295), .C(n297), .D(n309), .E(n299), .F(
        n310), .Z(n307) );
  GTECH_NOT U304 ( .A(n311), .Z(N148) );
  GTECH_AOI222 U305 ( .A(n312), .B(n295), .C(n297), .D(n313), .E(n299), .F(
        n314), .Z(n311) );
  GTECH_NOT U306 ( .A(n315), .Z(N147) );
  GTECH_AOI222 U307 ( .A(n316), .B(n295), .C(n297), .D(n317), .E(n299), .F(
        n318), .Z(n315) );
  GTECH_NOT U308 ( .A(n319), .Z(N146) );
  GTECH_AOI222 U309 ( .A(n320), .B(n295), .C(n297), .D(n321), .E(n299), .F(
        n322), .Z(n319) );
  GTECH_NOT U310 ( .A(n323), .Z(N145) );
  GTECH_AOI222 U311 ( .A(n324), .B(n295), .C(n297), .D(n325), .E(n299), .F(
        n326), .Z(n323) );
  GTECH_NOT U312 ( .A(n327), .Z(N144) );
  GTECH_AOI222 U313 ( .A(n328), .B(n295), .C(n297), .D(n329), .E(n299), .F(
        n330), .Z(n327) );
  GTECH_NOT U314 ( .A(n331), .Z(N143) );
  GTECH_AOI222 U315 ( .A(n332), .B(n295), .C(n297), .D(n333), .E(n299), .F(
        n334), .Z(n331) );
  GTECH_NOT U316 ( .A(n335), .Z(N142) );
  GTECH_AOI222 U317 ( .A(n336), .B(n295), .C(n297), .D(n337), .E(n299), .F(
        n338), .Z(n335) );
  GTECH_NOT U318 ( .A(n339), .Z(N141) );
  GTECH_AOI222 U319 ( .A(n340), .B(n295), .C(n297), .D(n341), .E(n299), .F(
        n342), .Z(n339) );
  GTECH_NOT U320 ( .A(n343), .Z(N140) );
  GTECH_AOI222 U321 ( .A(n344), .B(n295), .C(n297), .D(n345), .E(n299), .F(
        n346), .Z(n343) );
  GTECH_NOT U322 ( .A(n347), .Z(N14) );
  GTECH_NAND2 U323 ( .A(n286), .B(n249), .Z(n347) );
  GTECH_NOT U324 ( .A(n348), .Z(N139) );
  GTECH_AOI222 U325 ( .A(n349), .B(n295), .C(n297), .D(n350), .E(n299), .F(
        n351), .Z(n348) );
  GTECH_NOT U326 ( .A(n352), .Z(N138) );
  GTECH_AOI222 U327 ( .A(n353), .B(n295), .C(n297), .D(n354), .E(n299), .F(
        n355), .Z(n352) );
  GTECH_NOT U328 ( .A(n356), .Z(N137) );
  GTECH_AOI222 U329 ( .A(n357), .B(n295), .C(n297), .D(n358), .E(n299), .F(
        n359), .Z(n356) );
  GTECH_NOT U330 ( .A(n360), .Z(N136) );
  GTECH_AOI222 U331 ( .A(n295), .B(n269), .C(n297), .D(n271), .E(n299), .F(
        n273), .Z(n360) );
  GTECH_NOT U332 ( .A(n361), .Z(n273) );
  GTECH_XOR2 U333 ( .A(n362), .B(n363), .Z(n361) );
  GTECH_NOT U334 ( .A(n364), .Z(n363) );
  GTECH_NOT U335 ( .A(n365), .Z(n297) );
  GTECH_NOT U336 ( .A(n366), .Z(n269) );
  GTECH_XOR2 U337 ( .A(n362), .B(n367), .Z(n366) );
  GTECH_NOT U338 ( .A(n368), .Z(n367) );
  GTECH_XOR2 U339 ( .A(n271), .B(n251), .Z(n362) );
  GTECH_OAI21 U340 ( .A(n12), .B(n365), .C(n369), .Z(N135) );
  GTECH_OAI21 U341 ( .A(n299), .B(n295), .C(n277), .Z(n369) );
  GTECH_OAI21 U342 ( .A(n12), .B(n370), .C(n364), .Z(n277) );
  GTECH_NOT U343 ( .A(n371), .Z(n295) );
  GTECH_NAND3 U344 ( .A(n28), .B(n372), .C(N155), .Z(n371) );
  GTECH_NOT U345 ( .A(n373), .Z(n299) );
  GTECH_NAND3 U346 ( .A(n10), .B(n374), .C(N155), .Z(n373) );
  GTECH_NAND2 U347 ( .A(n375), .B(N155), .Z(n365) );
  GTECH_XOR2 U348 ( .A(n372), .B(n28), .Z(n375) );
  GTECH_AND2 U349 ( .A(N155), .B(n376), .Z(N134) );
  GTECH_NOT U350 ( .A(n13), .Z(n376) );
  GTECH_AND2 U351 ( .A(N155), .B(n377), .Z(N133) );
  GTECH_NOT U352 ( .A(n14), .Z(n377) );
  GTECH_AND2 U353 ( .A(N155), .B(n378), .Z(N132) );
  GTECH_NOT U354 ( .A(n15), .Z(n378) );
  GTECH_AND2 U355 ( .A(N155), .B(n379), .Z(N131) );
  GTECH_NOT U356 ( .A(n16), .Z(n379) );
  GTECH_AND2 U357 ( .A(N155), .B(n380), .Z(N130) );
  GTECH_NOT U358 ( .A(n17), .Z(n380) );
  GTECH_AND2 U359 ( .A(N155), .B(n381), .Z(N129) );
  GTECH_NOT U360 ( .A(n18), .Z(n381) );
  GTECH_AND2 U361 ( .A(N155), .B(n382), .Z(N128) );
  GTECH_NOT U362 ( .A(n19), .Z(n382) );
  GTECH_AND2 U363 ( .A(N155), .B(n383), .Z(N127) );
  GTECH_NOT U364 ( .A(n20), .Z(n383) );
  GTECH_AND2 U365 ( .A(N155), .B(n384), .Z(N126) );
  GTECH_NOT U366 ( .A(n21), .Z(n384) );
  GTECH_AND2 U367 ( .A(N155), .B(n385), .Z(N125) );
  GTECH_NOT U368 ( .A(n22), .Z(n385) );
  GTECH_AND2 U369 ( .A(N155), .B(n386), .Z(N124) );
  GTECH_NOT U370 ( .A(n23), .Z(n386) );
  GTECH_AND2 U371 ( .A(N155), .B(n387), .Z(N123) );
  GTECH_NOT U372 ( .A(n24), .Z(n387) );
  GTECH_AND2 U373 ( .A(N155), .B(n388), .Z(N122) );
  GTECH_NOT U374 ( .A(n25), .Z(n388) );
  GTECH_AND2 U375 ( .A(N155), .B(n389), .Z(N121) );
  GTECH_NOT U376 ( .A(n26), .Z(n389) );
  GTECH_AND2 U377 ( .A(N155), .B(n390), .Z(N120) );
  GTECH_NOT U378 ( .A(n27), .Z(n390) );
  GTECH_NOT U379 ( .A(n301), .Z(N155) );
  GTECH_NAND5 U380 ( .A(n391), .B(n6), .C(n9), .D(n8), .E(n7), .Z(n301) );
  GTECH_NOR2 U381 ( .A(n249), .B(Rst), .Z(n391) );
  GTECH_NOT U382 ( .A(n392), .Z(N116) );
  GTECH_AOI222 U383 ( .A(n270), .B(n298), .C(n272), .D(n300), .E(n296), .F(
        n268), .Z(n392) );
  GTECH_XOR2 U384 ( .A(n393), .B(n394), .Z(n296) );
  GTECH_ADD_ABC U385 ( .A(n31), .B(n265), .C(n395), .COUT(n394) );
  GTECH_XOR2 U386 ( .A(n396), .B(n393), .Z(n300) );
  GTECH_XOR2 U387 ( .A(A[16]), .B(n30), .Z(n393) );
  GTECH_OAI21 U388 ( .A(n397), .B(n31), .C(n398), .Z(n396) );
  GTECH_OAI21 U389 ( .A(n265), .B(n304), .C(n399), .Z(n398) );
  GTECH_NOT U390 ( .A(n30), .Z(n298) );
  GTECH_NAND2 U391 ( .A(n281), .B(n400), .Z(N115) );
  GTECH_NOT U392 ( .A(N41), .Z(n400) );
  GTECH_NAND2 U393 ( .A(n288), .B(n282), .Z(N41) );
  GTECH_NAND2 U394 ( .A(Ld), .B(n288), .Z(n282) );
  GTECH_NOT U395 ( .A(n401), .Z(N113) );
  GTECH_AOI222 U396 ( .A(n270), .B(n304), .C(n272), .D(n305), .E(n303), .F(
        n268), .Z(n401) );
  GTECH_XOR2 U397 ( .A(n402), .B(n395), .Z(n303) );
  GTECH_ADD_ABC U398 ( .A(n32), .B(n264), .C(n403), .COUT(n395) );
  GTECH_NOT U399 ( .A(n404), .Z(n305) );
  GTECH_XOR2 U400 ( .A(n402), .B(n405), .Z(n404) );
  GTECH_NOT U401 ( .A(n399), .Z(n405) );
  GTECH_OAI21 U402 ( .A(n32), .B(n406), .C(n407), .Z(n399) );
  GTECH_OAI21 U403 ( .A(n264), .B(n309), .C(n408), .Z(n407) );
  GTECH_XOR2 U404 ( .A(n397), .B(n31), .Z(n402) );
  GTECH_NOT U405 ( .A(n265), .Z(n397) );
  GTECH_NOT U406 ( .A(n31), .Z(n304) );
  GTECH_NOT U407 ( .A(n409), .Z(N112) );
  GTECH_AOI222 U408 ( .A(n270), .B(n309), .C(n272), .D(n310), .E(n308), .F(
        n268), .Z(n409) );
  GTECH_XOR2 U409 ( .A(n410), .B(n403), .Z(n308) );
  GTECH_ADD_ABC U410 ( .A(n33), .B(n263), .C(n411), .COUT(n403) );
  GTECH_NOT U411 ( .A(n412), .Z(n310) );
  GTECH_XOR2 U412 ( .A(n410), .B(n413), .Z(n412) );
  GTECH_NOT U413 ( .A(n408), .Z(n413) );
  GTECH_OAI21 U414 ( .A(n33), .B(n414), .C(n415), .Z(n408) );
  GTECH_OAI21 U415 ( .A(n263), .B(n313), .C(n416), .Z(n415) );
  GTECH_XOR2 U416 ( .A(n406), .B(n32), .Z(n410) );
  GTECH_NOT U417 ( .A(n264), .Z(n406) );
  GTECH_NOT U418 ( .A(n32), .Z(n309) );
  GTECH_NOT U419 ( .A(n417), .Z(N111) );
  GTECH_AOI222 U420 ( .A(n270), .B(n313), .C(n272), .D(n314), .E(n312), .F(
        n268), .Z(n417) );
  GTECH_XOR2 U421 ( .A(n418), .B(n411), .Z(n312) );
  GTECH_ADD_ABC U422 ( .A(n34), .B(n262), .C(n419), .COUT(n411) );
  GTECH_NOT U423 ( .A(n420), .Z(n314) );
  GTECH_XOR2 U424 ( .A(n418), .B(n421), .Z(n420) );
  GTECH_NOT U425 ( .A(n416), .Z(n421) );
  GTECH_OAI21 U426 ( .A(n34), .B(n422), .C(n423), .Z(n416) );
  GTECH_OAI21 U427 ( .A(n262), .B(n317), .C(n424), .Z(n423) );
  GTECH_XOR2 U428 ( .A(n414), .B(n33), .Z(n418) );
  GTECH_NOT U429 ( .A(n263), .Z(n414) );
  GTECH_NOT U430 ( .A(n33), .Z(n313) );
  GTECH_NOT U431 ( .A(n425), .Z(N110) );
  GTECH_AOI222 U432 ( .A(n270), .B(n317), .C(n272), .D(n318), .E(n316), .F(
        n268), .Z(n425) );
  GTECH_XOR2 U433 ( .A(n426), .B(n419), .Z(n316) );
  GTECH_ADD_ABC U434 ( .A(n35), .B(n261), .C(n427), .COUT(n419) );
  GTECH_NOT U435 ( .A(n428), .Z(n318) );
  GTECH_XOR2 U436 ( .A(n426), .B(n429), .Z(n428) );
  GTECH_NOT U437 ( .A(n424), .Z(n429) );
  GTECH_OAI21 U438 ( .A(n35), .B(n430), .C(n431), .Z(n424) );
  GTECH_OAI21 U439 ( .A(n261), .B(n321), .C(n432), .Z(n431) );
  GTECH_XOR2 U440 ( .A(n422), .B(n34), .Z(n426) );
  GTECH_NOT U441 ( .A(n262), .Z(n422) );
  GTECH_NOT U442 ( .A(n34), .Z(n317) );
  GTECH_NOT U443 ( .A(n433), .Z(N109) );
  GTECH_AOI222 U444 ( .A(n270), .B(n321), .C(n272), .D(n322), .E(n320), .F(
        n268), .Z(n433) );
  GTECH_XOR2 U445 ( .A(n434), .B(n427), .Z(n320) );
  GTECH_ADD_ABC U446 ( .A(n36), .B(n260), .C(n435), .COUT(n427) );
  GTECH_NOT U447 ( .A(n436), .Z(n322) );
  GTECH_XOR2 U448 ( .A(n434), .B(n437), .Z(n436) );
  GTECH_NOT U449 ( .A(n432), .Z(n437) );
  GTECH_OAI21 U450 ( .A(n36), .B(n438), .C(n439), .Z(n432) );
  GTECH_OAI21 U451 ( .A(n260), .B(n325), .C(n440), .Z(n439) );
  GTECH_XOR2 U452 ( .A(n430), .B(n35), .Z(n434) );
  GTECH_NOT U453 ( .A(n261), .Z(n430) );
  GTECH_NOT U454 ( .A(n35), .Z(n321) );
  GTECH_NOT U455 ( .A(n441), .Z(N108) );
  GTECH_AOI222 U456 ( .A(n270), .B(n325), .C(n272), .D(n326), .E(n324), .F(
        n268), .Z(n441) );
  GTECH_XOR2 U457 ( .A(n442), .B(n435), .Z(n324) );
  GTECH_ADD_ABC U458 ( .A(n37), .B(n259), .C(n443), .COUT(n435) );
  GTECH_NOT U459 ( .A(n444), .Z(n326) );
  GTECH_XOR2 U460 ( .A(n442), .B(n445), .Z(n444) );
  GTECH_NOT U461 ( .A(n440), .Z(n445) );
  GTECH_OAI21 U462 ( .A(n37), .B(n446), .C(n447), .Z(n440) );
  GTECH_OAI21 U463 ( .A(n259), .B(n329), .C(n448), .Z(n447) );
  GTECH_XOR2 U464 ( .A(n438), .B(n36), .Z(n442) );
  GTECH_NOT U465 ( .A(n260), .Z(n438) );
  GTECH_NOT U466 ( .A(n36), .Z(n325) );
  GTECH_NOT U467 ( .A(n449), .Z(N107) );
  GTECH_AOI222 U468 ( .A(n270), .B(n329), .C(n272), .D(n330), .E(n328), .F(
        n268), .Z(n449) );
  GTECH_XOR2 U469 ( .A(n450), .B(n443), .Z(n328) );
  GTECH_ADD_ABC U470 ( .A(n38), .B(n258), .C(n451), .COUT(n443) );
  GTECH_NOT U471 ( .A(n452), .Z(n330) );
  GTECH_XOR2 U472 ( .A(n450), .B(n453), .Z(n452) );
  GTECH_NOT U473 ( .A(n448), .Z(n453) );
  GTECH_OAI21 U474 ( .A(n38), .B(n454), .C(n455), .Z(n448) );
  GTECH_OAI21 U475 ( .A(n258), .B(n333), .C(n456), .Z(n455) );
  GTECH_XOR2 U476 ( .A(n446), .B(n37), .Z(n450) );
  GTECH_NOT U477 ( .A(n259), .Z(n446) );
  GTECH_NOT U478 ( .A(n37), .Z(n329) );
  GTECH_NOT U479 ( .A(n457), .Z(N106) );
  GTECH_AOI222 U480 ( .A(n270), .B(n333), .C(n272), .D(n334), .E(n332), .F(
        n268), .Z(n457) );
  GTECH_XOR2 U481 ( .A(n458), .B(n451), .Z(n332) );
  GTECH_ADD_ABC U482 ( .A(n39), .B(n257), .C(n459), .COUT(n451) );
  GTECH_NOT U483 ( .A(n460), .Z(n334) );
  GTECH_XOR2 U484 ( .A(n458), .B(n461), .Z(n460) );
  GTECH_NOT U485 ( .A(n456), .Z(n461) );
  GTECH_OAI21 U486 ( .A(n39), .B(n462), .C(n463), .Z(n456) );
  GTECH_OAI21 U487 ( .A(n257), .B(n337), .C(n464), .Z(n463) );
  GTECH_XOR2 U488 ( .A(n454), .B(n38), .Z(n458) );
  GTECH_NOT U489 ( .A(n258), .Z(n454) );
  GTECH_NOT U490 ( .A(n38), .Z(n333) );
  GTECH_NOT U491 ( .A(n465), .Z(N105) );
  GTECH_AOI222 U492 ( .A(n270), .B(n337), .C(n272), .D(n338), .E(n336), .F(
        n268), .Z(n465) );
  GTECH_XOR2 U493 ( .A(n466), .B(n459), .Z(n336) );
  GTECH_ADD_ABC U494 ( .A(n40), .B(n256), .C(n467), .COUT(n459) );
  GTECH_NOT U495 ( .A(n468), .Z(n338) );
  GTECH_XOR2 U496 ( .A(n466), .B(n469), .Z(n468) );
  GTECH_NOT U497 ( .A(n464), .Z(n469) );
  GTECH_OAI21 U498 ( .A(n40), .B(n470), .C(n471), .Z(n464) );
  GTECH_OAI21 U499 ( .A(n256), .B(n341), .C(n472), .Z(n471) );
  GTECH_XOR2 U500 ( .A(n462), .B(n39), .Z(n466) );
  GTECH_NOT U501 ( .A(n257), .Z(n462) );
  GTECH_NOT U502 ( .A(n39), .Z(n337) );
  GTECH_NOT U503 ( .A(n473), .Z(N104) );
  GTECH_AOI222 U504 ( .A(n270), .B(n341), .C(n272), .D(n342), .E(n340), .F(
        n268), .Z(n473) );
  GTECH_XOR2 U505 ( .A(n474), .B(n467), .Z(n340) );
  GTECH_ADD_ABC U506 ( .A(n41), .B(n255), .C(n475), .COUT(n467) );
  GTECH_NOT U507 ( .A(n476), .Z(n342) );
  GTECH_XOR2 U508 ( .A(n474), .B(n477), .Z(n476) );
  GTECH_NOT U509 ( .A(n472), .Z(n477) );
  GTECH_OAI21 U510 ( .A(n41), .B(n478), .C(n479), .Z(n472) );
  GTECH_OAI21 U511 ( .A(n255), .B(n345), .C(n480), .Z(n479) );
  GTECH_XOR2 U512 ( .A(n470), .B(n40), .Z(n474) );
  GTECH_NOT U513 ( .A(n256), .Z(n470) );
  GTECH_NOT U514 ( .A(n40), .Z(n341) );
  GTECH_NOT U515 ( .A(n481), .Z(N103) );
  GTECH_AOI222 U516 ( .A(n270), .B(n345), .C(n272), .D(n346), .E(n344), .F(
        n268), .Z(n481) );
  GTECH_XOR2 U517 ( .A(n482), .B(n475), .Z(n344) );
  GTECH_ADD_ABC U518 ( .A(n42), .B(n254), .C(n483), .COUT(n475) );
  GTECH_NOT U519 ( .A(n484), .Z(n346) );
  GTECH_XOR2 U520 ( .A(n482), .B(n485), .Z(n484) );
  GTECH_NOT U521 ( .A(n480), .Z(n485) );
  GTECH_OAI21 U522 ( .A(n42), .B(n486), .C(n487), .Z(n480) );
  GTECH_OAI21 U523 ( .A(n254), .B(n350), .C(n488), .Z(n487) );
  GTECH_XOR2 U524 ( .A(n478), .B(n41), .Z(n482) );
  GTECH_NOT U525 ( .A(n255), .Z(n478) );
  GTECH_NOT U526 ( .A(n41), .Z(n345) );
  GTECH_NOT U527 ( .A(n489), .Z(N102) );
  GTECH_AOI222 U528 ( .A(n270), .B(n350), .C(n272), .D(n351), .E(n349), .F(
        n268), .Z(n489) );
  GTECH_XOR2 U529 ( .A(n490), .B(n483), .Z(n349) );
  GTECH_ADD_ABC U530 ( .A(n43), .B(n253), .C(n491), .COUT(n483) );
  GTECH_NOT U531 ( .A(n492), .Z(n351) );
  GTECH_XOR2 U532 ( .A(n490), .B(n493), .Z(n492) );
  GTECH_NOT U533 ( .A(n488), .Z(n493) );
  GTECH_OAI21 U534 ( .A(n43), .B(n494), .C(n495), .Z(n488) );
  GTECH_OAI21 U535 ( .A(n253), .B(n354), .C(n496), .Z(n495) );
  GTECH_XOR2 U536 ( .A(n486), .B(n42), .Z(n490) );
  GTECH_NOT U537 ( .A(n254), .Z(n486) );
  GTECH_NOT U538 ( .A(n42), .Z(n350) );
  GTECH_NOT U539 ( .A(n497), .Z(N101) );
  GTECH_AOI222 U540 ( .A(n270), .B(n354), .C(n272), .D(n355), .E(n353), .F(
        n268), .Z(n497) );
  GTECH_XOR2 U541 ( .A(n498), .B(n491), .Z(n353) );
  GTECH_ADD_ABC U542 ( .A(n29), .B(n252), .C(n499), .COUT(n491) );
  GTECH_NOT U543 ( .A(n500), .Z(n355) );
  GTECH_XOR2 U544 ( .A(n498), .B(n501), .Z(n500) );
  GTECH_NOT U545 ( .A(n496), .Z(n501) );
  GTECH_OAI21 U546 ( .A(n29), .B(n502), .C(n503), .Z(n496) );
  GTECH_OAI21 U547 ( .A(n252), .B(n358), .C(n504), .Z(n503) );
  GTECH_XOR2 U548 ( .A(n494), .B(n43), .Z(n498) );
  GTECH_NOT U549 ( .A(n253), .Z(n494) );
  GTECH_NOT U550 ( .A(n43), .Z(n354) );
  GTECH_NOT U551 ( .A(n505), .Z(N100) );
  GTECH_AOI222 U552 ( .A(n357), .B(n268), .C(n270), .D(n358), .E(n272), .F(
        n359), .Z(n505) );
  GTECH_NOT U553 ( .A(n506), .Z(n359) );
  GTECH_XOR2 U554 ( .A(n507), .B(n508), .Z(n506) );
  GTECH_NOT U555 ( .A(n504), .Z(n508) );
  GTECH_OAI21 U556 ( .A(n11), .B(n509), .C(n510), .Z(n504) );
  GTECH_OAI21 U557 ( .A(n251), .B(n271), .C(n364), .Z(n510) );
  GTECH_NAND2 U558 ( .A(n12), .B(n370), .Z(n364) );
  GTECH_NOT U559 ( .A(n11), .Z(n271) );
  GTECH_NOT U560 ( .A(n251), .Z(n509) );
  GTECH_NOT U561 ( .A(n280), .Z(n272) );
  GTECH_NAND2 U562 ( .A(N82), .B(n10), .Z(n280) );
  GTECH_NOT U563 ( .A(n511), .Z(N82) );
  GTECH_NOT U564 ( .A(n29), .Z(n358) );
  GTECH_NOT U565 ( .A(n512), .Z(n270) );
  GTECH_MUX2 U566 ( .A(n511), .B(n513), .S(n10), .Z(n512) );
  GTECH_NAND2 U567 ( .A(n28), .B(n286), .Z(n513) );
  GTECH_NAND2 U568 ( .A(n286), .B(n374), .Z(n511) );
  GTECH_NOT U569 ( .A(n28), .Z(n374) );
  GTECH_NOT U570 ( .A(n279), .Z(n268) );
  GTECH_NAND3 U571 ( .A(n286), .B(n372), .C(n28), .Z(n279) );
  GTECH_NOT U572 ( .A(n10), .Z(n372) );
  GTECH_NOT U573 ( .A(n281), .Z(n286) );
  GTECH_OAI21 U574 ( .A(n284), .B(n285), .C(n514), .Z(n281) );
  GTECH_AND2 U575 ( .A(n287), .B(n288), .Z(n514) );
  GTECH_NOT U576 ( .A(Rst), .Z(n288) );
  GTECH_NOT U577 ( .A(Ld), .Z(n287) );
  GTECH_NOT U578 ( .A(n9), .Z(n285) );
  GTECH_NAND2 U579 ( .A(n8), .B(n290), .Z(n284) );
  GTECH_NOT U580 ( .A(n293), .Z(n290) );
  GTECH_NAND2 U581 ( .A(n7), .B(n292), .Z(n293) );
  GTECH_NOT U582 ( .A(n515), .Z(n292) );
  GTECH_NAND2 U583 ( .A(n6), .B(n249), .Z(n515) );
  GTECH_XOR2 U584 ( .A(n507), .B(n499), .Z(n357) );
  GTECH_ADD_ABC U585 ( .A(n251), .B(n11), .C(n368), .COUT(n499) );
  GTECH_NAND2 U586 ( .A(n275), .B(n370), .Z(n368) );
  GTECH_NOT U587 ( .A(n250), .Z(n370) );
  GTECH_NOT U588 ( .A(n12), .Z(n275) );
  GTECH_XOR2 U589 ( .A(n502), .B(n29), .Z(n507) );
  GTECH_NOT U590 ( .A(n252), .Z(n502) );
endmodule

