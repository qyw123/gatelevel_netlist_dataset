
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369;

  GTECH_MUX2 U131 ( .A(n270), .B(n271), .S(n272), .Z(sum[9]) );
  GTECH_XOR2 U132 ( .A(n273), .B(n274), .Z(n271) );
  GTECH_XOR2 U133 ( .A(n274), .B(n275), .Z(n270) );
  GTECH_AO21 U134 ( .A(a[9]), .B(b[9]), .C(n276), .Z(n274) );
  GTECH_XOR2 U135 ( .A(n272), .B(n277), .Z(sum[8]) );
  GTECH_MUX2 U136 ( .A(n278), .B(n279), .S(n280), .Z(sum[7]) );
  GTECH_XOR2 U137 ( .A(n281), .B(n282), .Z(n279) );
  GTECH_XNOR2 U138 ( .A(n281), .B(n283), .Z(n278) );
  GTECH_AOI21 U139 ( .A(n284), .B(n285), .C(n286), .Z(n283) );
  GTECH_XOR2 U140 ( .A(a[7]), .B(b[7]), .Z(n281) );
  GTECH_MUX2 U141 ( .A(n287), .B(n288), .S(n280), .Z(sum[6]) );
  GTECH_XNOR2 U142 ( .A(n289), .B(n290), .Z(n288) );
  GTECH_XNOR2 U143 ( .A(n285), .B(n289), .Z(n287) );
  GTECH_OR_NOT U144 ( .A(n286), .B(n284), .Z(n289) );
  GTECH_AO21 U145 ( .A(n291), .B(n292), .C(n293), .Z(n285) );
  GTECH_MUX2 U146 ( .A(n294), .B(n295), .S(n296), .Z(sum[5]) );
  GTECH_AND_NOT U147 ( .A(n291), .B(n293), .Z(n296) );
  GTECH_OAI21 U148 ( .A(n292), .B(n280), .C(n297), .Z(n295) );
  GTECH_AO21 U149 ( .A(n297), .B(n280), .C(n292), .Z(n294) );
  GTECH_XOR2 U150 ( .A(n280), .B(n298), .Z(sum[4]) );
  GTECH_MUX2 U151 ( .A(n299), .B(n300), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U152 ( .A(n301), .B(n302), .Z(n300) );
  GTECH_XNOR2 U153 ( .A(n301), .B(n303), .Z(n299) );
  GTECH_AOI21 U154 ( .A(n304), .B(n305), .C(n306), .Z(n303) );
  GTECH_XOR2 U155 ( .A(a[3]), .B(b[3]), .Z(n301) );
  GTECH_MUX2 U156 ( .A(n307), .B(n308), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U157 ( .A(n309), .B(n310), .Z(n308) );
  GTECH_XNOR2 U158 ( .A(n305), .B(n309), .Z(n307) );
  GTECH_OR_NOT U159 ( .A(n306), .B(n304), .Z(n309) );
  GTECH_OAI21 U160 ( .A(n311), .B(n312), .C(n313), .Z(n305) );
  GTECH_MUX2 U161 ( .A(n314), .B(n315), .S(n316), .Z(sum[1]) );
  GTECH_AND_NOT U162 ( .A(n313), .B(n311), .Z(n316) );
  GTECH_OAI21 U163 ( .A(cin), .B(n317), .C(n318), .Z(n315) );
  GTECH_AO21 U164 ( .A(n318), .B(cin), .C(n317), .Z(n314) );
  GTECH_NOT U165 ( .A(n312), .Z(n317) );
  GTECH_NAND2 U166 ( .A(a[0]), .B(b[0]), .Z(n312) );
  GTECH_MUX2 U167 ( .A(n319), .B(n320), .S(n321), .Z(sum[15]) );
  GTECH_XOR2 U168 ( .A(n322), .B(n323), .Z(n320) );
  GTECH_OA21 U169 ( .A(a[14]), .B(n324), .C(n325), .Z(n322) );
  GTECH_AO21 U170 ( .A(n324), .B(a[14]), .C(b[14]), .Z(n325) );
  GTECH_XNOR2 U171 ( .A(n323), .B(n326), .Z(n319) );
  GTECH_XOR2 U172 ( .A(n327), .B(n328), .Z(n323) );
  GTECH_MUX2 U173 ( .A(n329), .B(n330), .S(n321), .Z(sum[14]) );
  GTECH_XOR2 U174 ( .A(n331), .B(n324), .Z(n330) );
  GTECH_OAI2N2 U175 ( .A(n332), .B(n333), .C(a[13]), .D(b[13]), .Z(n324) );
  GTECH_XOR2 U176 ( .A(n331), .B(n334), .Z(n329) );
  GTECH_XOR2 U177 ( .A(a[14]), .B(b[14]), .Z(n331) );
  GTECH_MUX2 U178 ( .A(n335), .B(n336), .S(n321), .Z(sum[13]) );
  GTECH_XOR2 U179 ( .A(n333), .B(n337), .Z(n336) );
  GTECH_XOR2 U180 ( .A(n338), .B(n337), .Z(n335) );
  GTECH_AO21 U181 ( .A(a[13]), .B(b[13]), .C(n332), .Z(n337) );
  GTECH_NAND2 U182 ( .A(n339), .B(n340), .Z(sum[12]) );
  GTECH_AO21 U183 ( .A(n333), .B(n341), .C(n321), .Z(n339) );
  GTECH_MUX2 U184 ( .A(n342), .B(n343), .S(n272), .Z(sum[11]) );
  GTECH_XOR2 U185 ( .A(n344), .B(n345), .Z(n343) );
  GTECH_XNOR2 U186 ( .A(n344), .B(n346), .Z(n342) );
  GTECH_AOI21 U187 ( .A(n347), .B(n348), .C(n349), .Z(n346) );
  GTECH_XOR2 U188 ( .A(a[11]), .B(b[11]), .Z(n344) );
  GTECH_MUX2 U189 ( .A(n350), .B(n351), .S(n272), .Z(sum[10]) );
  GTECH_XNOR2 U190 ( .A(n352), .B(n353), .Z(n351) );
  GTECH_XNOR2 U191 ( .A(n348), .B(n353), .Z(n350) );
  GTECH_OR_NOT U192 ( .A(n349), .B(n347), .Z(n353) );
  GTECH_OAI2N2 U193 ( .A(n276), .B(n275), .C(a[9]), .D(b[9]), .Z(n348) );
  GTECH_XOR2 U194 ( .A(cin), .B(n354), .Z(sum[0]) );
  GTECH_OAI21 U195 ( .A(n355), .B(n321), .C(n340), .Z(cout) );
  GTECH_NAND3 U196 ( .A(n341), .B(n333), .C(n321), .Z(n340) );
  GTECH_NAND2 U197 ( .A(a[12]), .B(b[12]), .Z(n333) );
  GTECH_NOT U198 ( .A(n356), .Z(n321) );
  GTECH_MUX2 U199 ( .A(n277), .B(n357), .S(n272), .Z(n356) );
  GTECH_MUX2 U200 ( .A(n298), .B(n358), .S(n280), .Z(n272) );
  GTECH_MUX2 U201 ( .A(n354), .B(n359), .S(cin), .Z(n280) );
  GTECH_OA21 U202 ( .A(a[3]), .B(n302), .C(n360), .Z(n359) );
  GTECH_AO21 U203 ( .A(n302), .B(a[3]), .C(b[3]), .Z(n360) );
  GTECH_AO21 U204 ( .A(n310), .B(n304), .C(n306), .Z(n302) );
  GTECH_AND2 U205 ( .A(a[2]), .B(b[2]), .Z(n306) );
  GTECH_OR2 U206 ( .A(a[2]), .B(b[2]), .Z(n304) );
  GTECH_OAI21 U207 ( .A(n361), .B(n311), .C(n313), .Z(n310) );
  GTECH_NAND2 U208 ( .A(b[1]), .B(a[1]), .Z(n313) );
  GTECH_AND_NOT U209 ( .A(n362), .B(a[1]), .Z(n311) );
  GTECH_NOT U210 ( .A(b[1]), .Z(n362) );
  GTECH_NOT U211 ( .A(n318), .Z(n361) );
  GTECH_OR2 U212 ( .A(b[0]), .B(a[0]), .Z(n318) );
  GTECH_XOR2 U213 ( .A(a[0]), .B(b[0]), .Z(n354) );
  GTECH_OA21 U214 ( .A(a[7]), .B(n282), .C(n363), .Z(n358) );
  GTECH_AO21 U215 ( .A(n282), .B(a[7]), .C(b[7]), .Z(n363) );
  GTECH_AO21 U216 ( .A(n290), .B(n284), .C(n286), .Z(n282) );
  GTECH_AND2 U217 ( .A(a[6]), .B(b[6]), .Z(n286) );
  GTECH_OR2 U218 ( .A(a[6]), .B(b[6]), .Z(n284) );
  GTECH_AO21 U219 ( .A(n297), .B(n291), .C(n293), .Z(n290) );
  GTECH_AND2 U220 ( .A(a[5]), .B(b[5]), .Z(n293) );
  GTECH_OR2 U221 ( .A(b[5]), .B(a[5]), .Z(n291) );
  GTECH_AND_NOT U222 ( .A(n297), .B(n292), .Z(n298) );
  GTECH_AND2 U223 ( .A(b[4]), .B(a[4]), .Z(n292) );
  GTECH_OR2 U224 ( .A(a[4]), .B(b[4]), .Z(n297) );
  GTECH_OA21 U225 ( .A(a[11]), .B(n345), .C(n364), .Z(n357) );
  GTECH_AO21 U226 ( .A(n345), .B(a[11]), .C(b[11]), .Z(n364) );
  GTECH_AO21 U227 ( .A(n352), .B(n347), .C(n349), .Z(n345) );
  GTECH_AND2 U228 ( .A(a[10]), .B(b[10]), .Z(n349) );
  GTECH_OR2 U229 ( .A(a[10]), .B(b[10]), .Z(n347) );
  GTECH_OAI2N2 U230 ( .A(n276), .B(n273), .C(a[9]), .D(b[9]), .Z(n352) );
  GTECH_NOT U231 ( .A(n365), .Z(n273) );
  GTECH_NOT U232 ( .A(n366), .Z(n276) );
  GTECH_OR2 U233 ( .A(a[9]), .B(b[9]), .Z(n366) );
  GTECH_AND2 U234 ( .A(n275), .B(n365), .Z(n277) );
  GTECH_OR2 U235 ( .A(b[8]), .B(a[8]), .Z(n365) );
  GTECH_NAND2 U236 ( .A(a[8]), .B(b[8]), .Z(n275) );
  GTECH_OA21 U237 ( .A(n326), .B(n327), .C(n367), .Z(n355) );
  GTECH_AO21 U238 ( .A(n327), .B(n326), .C(n328), .Z(n367) );
  GTECH_NOT U239 ( .A(b[15]), .Z(n328) );
  GTECH_NOT U240 ( .A(a[15]), .Z(n327) );
  GTECH_AOI21 U241 ( .A(n334), .B(a[14]), .C(n368), .Z(n326) );
  GTECH_OA21 U242 ( .A(a[14]), .B(n334), .C(b[14]), .Z(n368) );
  GTECH_OAI2N2 U243 ( .A(n332), .B(n338), .C(a[13]), .D(b[13]), .Z(n334) );
  GTECH_NOT U244 ( .A(n341), .Z(n338) );
  GTECH_OR2 U245 ( .A(b[12]), .B(a[12]), .Z(n341) );
  GTECH_AND_NOT U246 ( .A(n369), .B(a[13]), .Z(n332) );
  GTECH_NOT U247 ( .A(b[13]), .Z(n369) );
endmodule

