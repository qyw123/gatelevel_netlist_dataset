
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_OR_NOT U83 ( .A(n97), .B(n93), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n98), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n98) );
  GTECH_OAI21 U86 ( .A(n99), .B(n100), .C(n101), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  GTECH_NOT U88 ( .A(n103), .Z(n99) );
  GTECH_OR_NOT U89 ( .A(n105), .B(I_b[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n106), .Z(n84) );
  GTECH_OR_NOT U91 ( .A(n107), .B(n108), .Z(n106) );
  GTECH_XOR2 U92 ( .A(n109), .B(n108), .Z(N153) );
  GTECH_NOT U93 ( .A(n110), .Z(n108) );
  GTECH_XOR3 U94 ( .A(n97), .B(n93), .C(n95), .Z(n110) );
  GTECH_XOR3 U95 ( .A(n102), .B(n104), .C(n103), .Z(n95) );
  GTECH_OAI21 U96 ( .A(n111), .B(n112), .C(n113), .Z(n103) );
  GTECH_OAI21 U97 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_NOT U98 ( .A(n115), .Z(n111) );
  GTECH_NOT U99 ( .A(n117), .Z(n104) );
  GTECH_OR_NOT U100 ( .A(n118), .B(I_b[7]), .Z(n117) );
  GTECH_NOT U101 ( .A(n100), .Z(n102) );
  GTECH_OR_NOT U102 ( .A(n119), .B(I_a[7]), .Z(n100) );
  GTECH_ADD_ABC U103 ( .A(n120), .B(n121), .C(n122), .COUT(n93) );
  GTECH_NOT U104 ( .A(n123), .Z(n122) );
  GTECH_XOR2 U105 ( .A(n124), .B(n125), .Z(n121) );
  GTECH_AND2 U106 ( .A(I_a[7]), .B(I_b[5]), .Z(n125) );
  GTECH_NOT U107 ( .A(n94), .Z(n97) );
  GTECH_OR_NOT U108 ( .A(n124), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U109 ( .A(n107), .Z(n109) );
  GTECH_OR_NOT U110 ( .A(n126), .B(n127), .Z(n107) );
  GTECH_XOR2 U111 ( .A(n126), .B(n128), .Z(N152) );
  GTECH_NOT U112 ( .A(n127), .Z(n128) );
  GTECH_XOR4 U113 ( .A(n129), .B(n124), .C(n120), .D(n123), .Z(n127) );
  GTECH_XOR3 U114 ( .A(n114), .B(n116), .C(n115), .Z(n123) );
  GTECH_OAI21 U115 ( .A(n130), .B(n131), .C(n132), .Z(n115) );
  GTECH_OAI21 U116 ( .A(n133), .B(n134), .C(n135), .Z(n132) );
  GTECH_NOT U117 ( .A(n134), .Z(n130) );
  GTECH_NOT U118 ( .A(n136), .Z(n116) );
  GTECH_OR_NOT U119 ( .A(n137), .B(I_b[7]), .Z(n136) );
  GTECH_NOT U120 ( .A(n112), .Z(n114) );
  GTECH_OR_NOT U121 ( .A(n118), .B(I_b[6]), .Z(n112) );
  GTECH_NOT U122 ( .A(I_a[6]), .Z(n118) );
  GTECH_ADD_ABC U123 ( .A(n138), .B(n139), .C(n140), .COUT(n120) );
  GTECH_NOT U124 ( .A(n141), .Z(n140) );
  GTECH_XOR3 U125 ( .A(n142), .B(n143), .C(n144), .Z(n139) );
  GTECH_OA21 U126 ( .A(n144), .B(n145), .C(n146), .Z(n124) );
  GTECH_OAI21 U127 ( .A(n142), .B(n147), .C(n143), .Z(n146) );
  GTECH_NOT U128 ( .A(n145), .Z(n142) );
  GTECH_NOT U129 ( .A(n147), .Z(n144) );
  GTECH_AND2 U130 ( .A(I_b[5]), .B(I_a[7]), .Z(n129) );
  GTECH_ADD_ABC U131 ( .A(n148), .B(n149), .C(n150), .COUT(n126) );
  GTECH_NOT U132 ( .A(n151), .Z(n150) );
  GTECH_OA22 U133 ( .A(n152), .B(n105), .C(n153), .D(n154), .Z(n149) );
  GTECH_OA21 U134 ( .A(n155), .B(n156), .C(n157), .Z(n148) );
  GTECH_XOR3 U135 ( .A(n158), .B(n151), .C(n159), .Z(N151) );
  GTECH_OA21 U136 ( .A(n155), .B(n156), .C(n157), .Z(n159) );
  GTECH_OAI21 U137 ( .A(n160), .B(n161), .C(n162), .Z(n157) );
  GTECH_XOR2 U138 ( .A(n163), .B(n138), .Z(n151) );
  GTECH_ADD_ABC U139 ( .A(n164), .B(n165), .C(n166), .COUT(n138) );
  GTECH_NOT U140 ( .A(n167), .Z(n166) );
  GTECH_XOR3 U141 ( .A(n168), .B(n169), .C(n170), .Z(n165) );
  GTECH_XOR4 U142 ( .A(n143), .B(n147), .C(n145), .D(n141), .Z(n163) );
  GTECH_XOR3 U143 ( .A(n133), .B(n135), .C(n134), .Z(n141) );
  GTECH_OAI21 U144 ( .A(n171), .B(n172), .C(n173), .Z(n134) );
  GTECH_OAI21 U145 ( .A(n174), .B(n175), .C(n176), .Z(n173) );
  GTECH_NOT U146 ( .A(n175), .Z(n171) );
  GTECH_NOT U147 ( .A(n177), .Z(n135) );
  GTECH_OR_NOT U148 ( .A(n178), .B(I_b[7]), .Z(n177) );
  GTECH_NOT U149 ( .A(n131), .Z(n133) );
  GTECH_OR_NOT U150 ( .A(n137), .B(I_b[6]), .Z(n131) );
  GTECH_NOT U151 ( .A(I_a[5]), .Z(n137) );
  GTECH_OR_NOT U152 ( .A(n179), .B(I_a[7]), .Z(n145) );
  GTECH_OAI21 U153 ( .A(n170), .B(n180), .C(n181), .Z(n147) );
  GTECH_OAI21 U154 ( .A(n168), .B(n182), .C(n169), .Z(n181) );
  GTECH_NOT U155 ( .A(n180), .Z(n168) );
  GTECH_NOT U156 ( .A(n182), .Z(n170) );
  GTECH_NOT U157 ( .A(n183), .Z(n143) );
  GTECH_OR_NOT U158 ( .A(n184), .B(I_a[6]), .Z(n183) );
  GTECH_OA22 U159 ( .A(n152), .B(n105), .C(n153), .D(n154), .Z(n158) );
  GTECH_NOT U160 ( .A(n185), .Z(n154) );
  GTECH_NOT U161 ( .A(I_a[7]), .Z(n105) );
  GTECH_XOR3 U162 ( .A(n155), .B(n160), .C(n186), .Z(N150) );
  GTECH_NOT U163 ( .A(n162), .Z(n186) );
  GTECH_XOR2 U164 ( .A(n187), .B(n164), .Z(n162) );
  GTECH_ADD_ABC U165 ( .A(n188), .B(n189), .C(n190), .COUT(n164) );
  GTECH_NOT U166 ( .A(n191), .Z(n190) );
  GTECH_XOR3 U167 ( .A(n192), .B(n193), .C(n194), .Z(n189) );
  GTECH_XOR4 U168 ( .A(n169), .B(n182), .C(n180), .D(n167), .Z(n187) );
  GTECH_XOR3 U169 ( .A(n174), .B(n176), .C(n175), .Z(n167) );
  GTECH_OAI21 U170 ( .A(n195), .B(n196), .C(n197), .Z(n175) );
  GTECH_OAI21 U171 ( .A(n198), .B(n199), .C(n200), .Z(n197) );
  GTECH_NOT U172 ( .A(n199), .Z(n195) );
  GTECH_NOT U173 ( .A(n201), .Z(n176) );
  GTECH_OR_NOT U174 ( .A(n202), .B(I_b[7]), .Z(n201) );
  GTECH_NOT U175 ( .A(n172), .Z(n174) );
  GTECH_OR_NOT U176 ( .A(n178), .B(I_b[6]), .Z(n172) );
  GTECH_OR_NOT U177 ( .A(n179), .B(I_a[6]), .Z(n180) );
  GTECH_OAI21 U178 ( .A(n194), .B(n203), .C(n204), .Z(n182) );
  GTECH_OAI21 U179 ( .A(n192), .B(n205), .C(n193), .Z(n204) );
  GTECH_NOT U180 ( .A(n203), .Z(n192) );
  GTECH_NOT U181 ( .A(n205), .Z(n194) );
  GTECH_NOT U182 ( .A(n206), .Z(n169) );
  GTECH_OR_NOT U183 ( .A(n184), .B(I_a[5]), .Z(n206) );
  GTECH_NOT U184 ( .A(I_b[5]), .Z(n184) );
  GTECH_NOT U185 ( .A(n156), .Z(n160) );
  GTECH_XOR2 U186 ( .A(n185), .B(n153), .Z(n156) );
  GTECH_AOI2N2 U187 ( .A(n207), .B(n208), .C(n209), .D(n210), .Z(n153) );
  GTECH_OR_NOT U188 ( .A(n211), .B(n209), .Z(n208) );
  GTECH_XOR2 U189 ( .A(n212), .B(n152), .Z(n185) );
  GTECH_AND2 U190 ( .A(n213), .B(n214), .Z(n152) );
  GTECH_OR_NOT U191 ( .A(n215), .B(n216), .Z(n214) );
  GTECH_OAI21 U192 ( .A(n217), .B(n216), .C(n218), .Z(n213) );
  GTECH_OR_NOT U193 ( .A(n219), .B(I_a[7]), .Z(n212) );
  GTECH_NOT U194 ( .A(n161), .Z(n155) );
  GTECH_OAI2N2 U195 ( .A(n220), .B(n221), .C(n222), .D(n223), .Z(n161) );
  GTECH_OR_NOT U196 ( .A(n224), .B(n220), .Z(n223) );
  GTECH_XOR3 U197 ( .A(n220), .B(n224), .C(n225), .Z(N149) );
  GTECH_NOT U198 ( .A(n222), .Z(n225) );
  GTECH_XOR2 U199 ( .A(n226), .B(n188), .Z(n222) );
  GTECH_ADD_ABC U200 ( .A(n227), .B(n228), .C(n229), .COUT(n188) );
  GTECH_XOR3 U201 ( .A(n230), .B(n231), .C(n232), .Z(n228) );
  GTECH_OA21 U202 ( .A(n233), .B(n234), .C(n235), .Z(n227) );
  GTECH_XOR4 U203 ( .A(n193), .B(n205), .C(n203), .D(n191), .Z(n226) );
  GTECH_XOR3 U204 ( .A(n198), .B(n200), .C(n199), .Z(n191) );
  GTECH_OAI21 U205 ( .A(n236), .B(n237), .C(n238), .Z(n199) );
  GTECH_NOT U206 ( .A(n239), .Z(n200) );
  GTECH_OR_NOT U207 ( .A(n240), .B(I_b[7]), .Z(n239) );
  GTECH_NOT U208 ( .A(n196), .Z(n198) );
  GTECH_OR_NOT U209 ( .A(n202), .B(I_b[6]), .Z(n196) );
  GTECH_OR_NOT U210 ( .A(n179), .B(I_a[5]), .Z(n203) );
  GTECH_OAI21 U211 ( .A(n232), .B(n241), .C(n242), .Z(n205) );
  GTECH_OAI21 U212 ( .A(n230), .B(n243), .C(n231), .Z(n242) );
  GTECH_NOT U213 ( .A(n241), .Z(n230) );
  GTECH_NOT U214 ( .A(n243), .Z(n232) );
  GTECH_NOT U215 ( .A(n244), .Z(n193) );
  GTECH_OR_NOT U216 ( .A(n178), .B(I_b[5]), .Z(n244) );
  GTECH_NOT U217 ( .A(n221), .Z(n224) );
  GTECH_XOR3 U218 ( .A(n211), .B(n209), .C(n207), .Z(n221) );
  GTECH_XOR3 U219 ( .A(n217), .B(n218), .C(n216), .Z(n207) );
  GTECH_OAI21 U220 ( .A(n245), .B(n246), .C(n247), .Z(n216) );
  GTECH_OAI21 U221 ( .A(n248), .B(n249), .C(n250), .Z(n247) );
  GTECH_NOT U222 ( .A(n249), .Z(n245) );
  GTECH_NOT U223 ( .A(n251), .Z(n218) );
  GTECH_OR_NOT U224 ( .A(n219), .B(I_a[6]), .Z(n251) );
  GTECH_NOT U225 ( .A(n215), .Z(n217) );
  GTECH_OR_NOT U226 ( .A(n252), .B(I_a[7]), .Z(n215) );
  GTECH_ADD_ABC U227 ( .A(n253), .B(n254), .C(n255), .COUT(n209) );
  GTECH_XOR2 U228 ( .A(n256), .B(n257), .Z(n254) );
  GTECH_AND2 U229 ( .A(I_a[7]), .B(I_b[1]), .Z(n257) );
  GTECH_NOT U230 ( .A(n210), .Z(n211) );
  GTECH_OR_NOT U231 ( .A(n256), .B(I_a[7]), .Z(n210) );
  GTECH_ADD_ABC U232 ( .A(n258), .B(n259), .C(n260), .COUT(n220) );
  GTECH_XOR3 U233 ( .A(n253), .B(n261), .C(n255), .Z(n259) );
  GTECH_NOT U234 ( .A(n262), .Z(n255) );
  GTECH_XOR2 U235 ( .A(n258), .B(n263), .Z(N148) );
  GTECH_XOR4 U236 ( .A(n261), .B(n262), .C(n260), .D(n253), .Z(n263) );
  GTECH_ADD_ABC U237 ( .A(n264), .B(n265), .C(n266), .COUT(n253) );
  GTECH_XOR3 U238 ( .A(n267), .B(n268), .C(n269), .Z(n265) );
  GTECH_XOR2 U239 ( .A(n270), .B(n271), .Z(n260) );
  GTECH_OA21 U240 ( .A(n233), .B(n234), .C(n235), .Z(n271) );
  GTECH_OAI21 U241 ( .A(n272), .B(n273), .C(n274), .Z(n235) );
  GTECH_NOT U242 ( .A(n233), .Z(n273) );
  GTECH_XOR4 U243 ( .A(n231), .B(n243), .C(n241), .D(n229), .Z(n270) );
  GTECH_XOR3 U244 ( .A(n275), .B(n276), .C(n238), .Z(n229) );
  GTECH_OR3 U245 ( .A(n277), .B(n119), .C(n278), .Z(n238) );
  GTECH_NOT U246 ( .A(n237), .Z(n276) );
  GTECH_OR_NOT U247 ( .A(n277), .B(I_b[7]), .Z(n237) );
  GTECH_NOT U248 ( .A(n236), .Z(n275) );
  GTECH_OR_NOT U249 ( .A(n240), .B(I_b[6]), .Z(n236) );
  GTECH_OR_NOT U250 ( .A(n178), .B(I_b[4]), .Z(n241) );
  GTECH_OAI21 U251 ( .A(n279), .B(n280), .C(n281), .Z(n243) );
  GTECH_OAI21 U252 ( .A(n282), .B(n283), .C(n284), .Z(n281) );
  GTECH_NOT U253 ( .A(n283), .Z(n279) );
  GTECH_NOT U254 ( .A(n285), .Z(n231) );
  GTECH_OR_NOT U255 ( .A(n202), .B(I_b[5]), .Z(n285) );
  GTECH_XOR3 U256 ( .A(n248), .B(n250), .C(n249), .Z(n262) );
  GTECH_OAI21 U257 ( .A(n286), .B(n287), .C(n288), .Z(n249) );
  GTECH_OAI21 U258 ( .A(n289), .B(n290), .C(n291), .Z(n288) );
  GTECH_NOT U259 ( .A(n290), .Z(n286) );
  GTECH_NOT U260 ( .A(n292), .Z(n250) );
  GTECH_OR_NOT U261 ( .A(n219), .B(I_a[5]), .Z(n292) );
  GTECH_NOT U262 ( .A(I_b[3]), .Z(n219) );
  GTECH_NOT U263 ( .A(n246), .Z(n248) );
  GTECH_OR_NOT U264 ( .A(n252), .B(I_a[6]), .Z(n246) );
  GTECH_XOR2 U265 ( .A(n293), .B(n256), .Z(n261) );
  GTECH_OA21 U266 ( .A(n269), .B(n294), .C(n295), .Z(n256) );
  GTECH_OAI21 U267 ( .A(n267), .B(n296), .C(n268), .Z(n295) );
  GTECH_NOT U268 ( .A(n296), .Z(n269) );
  GTECH_AND2 U269 ( .A(I_b[1]), .B(I_a[7]), .Z(n293) );
  GTECH_ADD_ABC U270 ( .A(n297), .B(n298), .C(n299), .COUT(n258) );
  GTECH_NOT U271 ( .A(n300), .Z(n299) );
  GTECH_XOR3 U272 ( .A(n264), .B(n301), .C(n266), .Z(n298) );
  GTECH_NOT U273 ( .A(n302), .Z(n266) );
  GTECH_NOT U274 ( .A(n303), .Z(n301) );
  GTECH_XOR2 U275 ( .A(n304), .B(n297), .Z(N147) );
  GTECH_ADD_ABC U276 ( .A(n305), .B(n306), .C(n307), .COUT(n297) );
  GTECH_XOR3 U277 ( .A(n308), .B(n309), .C(n310), .Z(n306) );
  GTECH_OA21 U278 ( .A(n311), .B(n312), .C(n313), .Z(n305) );
  GTECH_XOR4 U279 ( .A(n302), .B(n264), .C(n303), .D(n300), .Z(n304) );
  GTECH_XOR3 U280 ( .A(n274), .B(n234), .C(n233), .Z(n300) );
  GTECH_XOR2 U281 ( .A(n314), .B(n278), .Z(n233) );
  GTECH_OR_NOT U282 ( .A(n315), .B(I_b[7]), .Z(n278) );
  GTECH_AND2 U283 ( .A(I_a[1]), .B(I_b[6]), .Z(n314) );
  GTECH_NOT U284 ( .A(n272), .Z(n234) );
  GTECH_XOR3 U285 ( .A(n282), .B(n284), .C(n283), .Z(n272) );
  GTECH_OAI21 U286 ( .A(n316), .B(n317), .C(n318), .Z(n283) );
  GTECH_NOT U287 ( .A(n319), .Z(n284) );
  GTECH_OR_NOT U288 ( .A(n240), .B(I_b[5]), .Z(n319) );
  GTECH_NOT U289 ( .A(n280), .Z(n282) );
  GTECH_OR_NOT U290 ( .A(n202), .B(I_b[4]), .Z(n280) );
  GTECH_NOT U291 ( .A(n320), .Z(n274) );
  GTECH_OR3 U292 ( .A(n321), .B(n315), .C(n119), .Z(n320) );
  GTECH_NOT U293 ( .A(I_b[6]), .Z(n119) );
  GTECH_XOR3 U294 ( .A(n267), .B(n268), .C(n296), .Z(n303) );
  GTECH_OAI21 U295 ( .A(n322), .B(n323), .C(n324), .Z(n296) );
  GTECH_OAI21 U296 ( .A(n325), .B(n326), .C(n327), .Z(n324) );
  GTECH_NOT U297 ( .A(n328), .Z(n268) );
  GTECH_OR_NOT U298 ( .A(n329), .B(I_a[6]), .Z(n328) );
  GTECH_NOT U299 ( .A(n294), .Z(n267) );
  GTECH_OR_NOT U300 ( .A(n330), .B(I_a[7]), .Z(n294) );
  GTECH_ADD_ABC U301 ( .A(n308), .B(n331), .C(n310), .COUT(n264) );
  GTECH_NOT U302 ( .A(n332), .Z(n310) );
  GTECH_XOR3 U303 ( .A(n325), .B(n327), .C(n322), .Z(n331) );
  GTECH_NOT U304 ( .A(n326), .Z(n322) );
  GTECH_XOR3 U305 ( .A(n289), .B(n291), .C(n290), .Z(n302) );
  GTECH_OAI21 U306 ( .A(n333), .B(n334), .C(n335), .Z(n290) );
  GTECH_OAI21 U307 ( .A(n336), .B(n337), .C(n338), .Z(n335) );
  GTECH_NOT U308 ( .A(n337), .Z(n333) );
  GTECH_NOT U309 ( .A(n339), .Z(n291) );
  GTECH_OR_NOT U310 ( .A(n178), .B(I_b[3]), .Z(n339) );
  GTECH_NOT U311 ( .A(n287), .Z(n289) );
  GTECH_OR_NOT U312 ( .A(n252), .B(I_a[5]), .Z(n287) );
  GTECH_XOR2 U313 ( .A(n340), .B(n341), .Z(N146) );
  GTECH_XOR4 U314 ( .A(n309), .B(n332), .C(n307), .D(n308), .Z(n341) );
  GTECH_ADD_ABC U315 ( .A(n342), .B(n343), .C(n344), .COUT(n308) );
  GTECH_NOT U316 ( .A(n345), .Z(n344) );
  GTECH_XOR3 U317 ( .A(n346), .B(n347), .C(n348), .Z(n343) );
  GTECH_XOR2 U318 ( .A(n321), .B(n349), .Z(n307) );
  GTECH_AND2 U319 ( .A(I_b[6]), .B(I_a[0]), .Z(n349) );
  GTECH_XOR3 U320 ( .A(n350), .B(n351), .C(n318), .Z(n321) );
  GTECH_OR3 U321 ( .A(n277), .B(n179), .C(n352), .Z(n318) );
  GTECH_NOT U322 ( .A(n317), .Z(n351) );
  GTECH_OR_NOT U323 ( .A(n277), .B(I_b[5]), .Z(n317) );
  GTECH_NOT U324 ( .A(n316), .Z(n350) );
  GTECH_OR_NOT U325 ( .A(n240), .B(I_b[4]), .Z(n316) );
  GTECH_XOR3 U326 ( .A(n336), .B(n338), .C(n337), .Z(n332) );
  GTECH_OAI21 U327 ( .A(n353), .B(n354), .C(n355), .Z(n337) );
  GTECH_OAI21 U328 ( .A(n356), .B(n357), .C(n358), .Z(n355) );
  GTECH_NOT U329 ( .A(n357), .Z(n353) );
  GTECH_NOT U330 ( .A(n359), .Z(n338) );
  GTECH_OR_NOT U331 ( .A(n202), .B(I_b[3]), .Z(n359) );
  GTECH_NOT U332 ( .A(n334), .Z(n336) );
  GTECH_OR_NOT U333 ( .A(n178), .B(I_b[2]), .Z(n334) );
  GTECH_NOT U334 ( .A(I_a[4]), .Z(n178) );
  GTECH_NOT U335 ( .A(n360), .Z(n309) );
  GTECH_XOR3 U336 ( .A(n325), .B(n327), .C(n326), .Z(n360) );
  GTECH_OAI21 U337 ( .A(n348), .B(n361), .C(n362), .Z(n326) );
  GTECH_OAI21 U338 ( .A(n346), .B(n363), .C(n347), .Z(n362) );
  GTECH_NOT U339 ( .A(n361), .Z(n346) );
  GTECH_NOT U340 ( .A(n363), .Z(n348) );
  GTECH_NOT U341 ( .A(n364), .Z(n327) );
  GTECH_OR_NOT U342 ( .A(n329), .B(I_a[5]), .Z(n364) );
  GTECH_NOT U343 ( .A(n323), .Z(n325) );
  GTECH_OR_NOT U344 ( .A(n330), .B(I_a[6]), .Z(n323) );
  GTECH_OA21 U345 ( .A(n311), .B(n312), .C(n313), .Z(n340) );
  GTECH_OAI21 U346 ( .A(n365), .B(n366), .C(n367), .Z(n313) );
  GTECH_NOT U347 ( .A(n311), .Z(n366) );
  GTECH_XOR3 U348 ( .A(n367), .B(n312), .C(n311), .Z(N145) );
  GTECH_XOR2 U349 ( .A(n368), .B(n352), .Z(n311) );
  GTECH_OR_NOT U350 ( .A(n315), .B(I_b[5]), .Z(n352) );
  GTECH_AND2 U351 ( .A(I_a[1]), .B(I_b[4]), .Z(n368) );
  GTECH_NOT U352 ( .A(n365), .Z(n312) );
  GTECH_XOR2 U353 ( .A(n369), .B(n342), .Z(n365) );
  GTECH_ADD_ABC U354 ( .A(n370), .B(n371), .C(n372), .COUT(n342) );
  GTECH_XOR3 U355 ( .A(n373), .B(n374), .C(n375), .Z(n371) );
  GTECH_OA21 U356 ( .A(n376), .B(n377), .C(n378), .Z(n370) );
  GTECH_XOR4 U357 ( .A(n347), .B(n363), .C(n361), .D(n345), .Z(n369) );
  GTECH_XOR3 U358 ( .A(n356), .B(n358), .C(n357), .Z(n345) );
  GTECH_OAI21 U359 ( .A(n379), .B(n380), .C(n381), .Z(n357) );
  GTECH_NOT U360 ( .A(n382), .Z(n358) );
  GTECH_OR_NOT U361 ( .A(n240), .B(I_b[3]), .Z(n382) );
  GTECH_NOT U362 ( .A(n354), .Z(n356) );
  GTECH_OR_NOT U363 ( .A(n202), .B(I_b[2]), .Z(n354) );
  GTECH_OR_NOT U364 ( .A(n330), .B(I_a[5]), .Z(n361) );
  GTECH_OAI21 U365 ( .A(n375), .B(n383), .C(n384), .Z(n363) );
  GTECH_OAI21 U366 ( .A(n373), .B(n385), .C(n374), .Z(n384) );
  GTECH_NOT U367 ( .A(n383), .Z(n373) );
  GTECH_NOT U368 ( .A(n385), .Z(n375) );
  GTECH_NOT U369 ( .A(n386), .Z(n347) );
  GTECH_OR_NOT U370 ( .A(n329), .B(I_a[4]), .Z(n386) );
  GTECH_NOT U371 ( .A(n387), .Z(n367) );
  GTECH_OR3 U372 ( .A(n388), .B(n315), .C(n179), .Z(n387) );
  GTECH_NOT U373 ( .A(I_b[4]), .Z(n179) );
  GTECH_XNOR2 U374 ( .A(n389), .B(n388), .Z(N144) );
  GTECH_XOR2 U375 ( .A(n390), .B(n391), .Z(n388) );
  GTECH_OA21 U376 ( .A(n376), .B(n377), .C(n378), .Z(n391) );
  GTECH_OAI21 U377 ( .A(n392), .B(n393), .C(n394), .Z(n378) );
  GTECH_NOT U378 ( .A(n376), .Z(n393) );
  GTECH_XOR4 U379 ( .A(n374), .B(n385), .C(n383), .D(n372), .Z(n390) );
  GTECH_XOR3 U380 ( .A(n395), .B(n396), .C(n381), .Z(n372) );
  GTECH_OR3 U381 ( .A(n277), .B(n252), .C(n397), .Z(n381) );
  GTECH_NOT U382 ( .A(n380), .Z(n396) );
  GTECH_OR_NOT U383 ( .A(n277), .B(I_b[3]), .Z(n380) );
  GTECH_NOT U384 ( .A(n379), .Z(n395) );
  GTECH_OR_NOT U385 ( .A(n240), .B(I_b[2]), .Z(n379) );
  GTECH_OR_NOT U386 ( .A(n330), .B(I_a[4]), .Z(n383) );
  GTECH_OAI21 U387 ( .A(n398), .B(n399), .C(n400), .Z(n385) );
  GTECH_OAI21 U388 ( .A(n401), .B(n402), .C(n403), .Z(n400) );
  GTECH_NOT U389 ( .A(n402), .Z(n398) );
  GTECH_NOT U390 ( .A(n404), .Z(n374) );
  GTECH_OR_NOT U391 ( .A(n329), .B(I_a[3]), .Z(n404) );
  GTECH_AND2 U392 ( .A(I_b[4]), .B(I_a[0]), .Z(n389) );
  GTECH_XOR3 U393 ( .A(n394), .B(n377), .C(n376), .Z(N143) );
  GTECH_XOR2 U394 ( .A(n405), .B(n397), .Z(n376) );
  GTECH_OR_NOT U395 ( .A(n315), .B(I_b[3]), .Z(n397) );
  GTECH_AND2 U396 ( .A(I_a[1]), .B(I_b[2]), .Z(n405) );
  GTECH_NOT U397 ( .A(n392), .Z(n377) );
  GTECH_XOR3 U398 ( .A(n401), .B(n403), .C(n402), .Z(n392) );
  GTECH_OAI21 U399 ( .A(n406), .B(n407), .C(n408), .Z(n402) );
  GTECH_NOT U400 ( .A(n409), .Z(n403) );
  GTECH_OR_NOT U401 ( .A(n240), .B(I_b[1]), .Z(n409) );
  GTECH_NOT U402 ( .A(n399), .Z(n401) );
  GTECH_OR_NOT U403 ( .A(n202), .B(I_b[0]), .Z(n399) );
  GTECH_NOT U404 ( .A(I_a[3]), .Z(n202) );
  GTECH_NOT U405 ( .A(n410), .Z(n394) );
  GTECH_OR3 U406 ( .A(n411), .B(n315), .C(n252), .Z(n410) );
  GTECH_NOT U407 ( .A(I_b[2]), .Z(n252) );
  GTECH_NOT U408 ( .A(I_a[0]), .Z(n315) );
  GTECH_XNOR2 U409 ( .A(n412), .B(n411), .Z(N142) );
  GTECH_XOR3 U410 ( .A(n413), .B(n414), .C(n408), .Z(n411) );
  GTECH_OR3 U411 ( .A(n330), .B(n415), .C(n277), .Z(n408) );
  GTECH_NOT U412 ( .A(I_a[1]), .Z(n277) );
  GTECH_NOT U413 ( .A(I_b[0]), .Z(n330) );
  GTECH_NOT U414 ( .A(n406), .Z(n414) );
  GTECH_OR_NOT U415 ( .A(n329), .B(I_a[1]), .Z(n406) );
  GTECH_NOT U416 ( .A(n407), .Z(n413) );
  GTECH_OR_NOT U417 ( .A(n240), .B(I_b[0]), .Z(n407) );
  GTECH_NOT U418 ( .A(I_a[2]), .Z(n240) );
  GTECH_AND2 U419 ( .A(I_b[2]), .B(I_a[0]), .Z(n412) );
  GTECH_XNOR2 U420 ( .A(n415), .B(n416), .Z(N141) );
  GTECH_AND2 U421 ( .A(I_a[1]), .B(I_b[0]), .Z(n416) );
  GTECH_OR_NOT U422 ( .A(n329), .B(I_a[0]), .Z(n415) );
  GTECH_NOT U423 ( .A(I_b[1]), .Z(n329) );
  GTECH_AND2 U424 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

