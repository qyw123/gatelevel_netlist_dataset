
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389;

  GTECH_MUX2 U136 ( .A(n275), .B(n276), .S(n277), .Z(sum[9]) );
  GTECH_XOR2 U137 ( .A(n278), .B(n279), .Z(n276) );
  GTECH_XOR2 U138 ( .A(n279), .B(n280), .Z(n275) );
  GTECH_AND_NOT U139 ( .A(n281), .B(n282), .Z(n279) );
  GTECH_XOR2 U140 ( .A(n283), .B(n284), .Z(sum[8]) );
  GTECH_MUX2 U141 ( .A(n285), .B(n286), .S(n287), .Z(sum[7]) );
  GTECH_XNOR2 U142 ( .A(n288), .B(n289), .Z(n286) );
  GTECH_OA21 U143 ( .A(n290), .B(n291), .C(n292), .Z(n289) );
  GTECH_XOR2 U144 ( .A(n288), .B(n293), .Z(n285) );
  GTECH_XOR2 U145 ( .A(a[7]), .B(b[7]), .Z(n288) );
  GTECH_MUX2 U146 ( .A(n294), .B(n295), .S(n287), .Z(sum[6]) );
  GTECH_XNOR2 U147 ( .A(n296), .B(n291), .Z(n295) );
  GTECH_AOI21 U148 ( .A(a[4]), .B(n297), .C(n298), .Z(n291) );
  GTECH_AND_NOT U149 ( .A(b[4]), .B(n299), .Z(n297) );
  GTECH_XNOR2 U150 ( .A(n296), .B(n300), .Z(n294) );
  GTECH_NOR2 U151 ( .A(n301), .B(n290), .Z(n296) );
  GTECH_XOR2 U152 ( .A(n302), .B(n303), .Z(sum[5]) );
  GTECH_AND_NOT U153 ( .A(n304), .B(n299), .Z(n303) );
  GTECH_ADD_ABC U154 ( .A(a[4]), .B(n305), .C(b[4]), .COUT(n302) );
  GTECH_MUX2 U155 ( .A(n306), .B(n307), .S(cin), .Z(n305) );
  GTECH_OAI21 U156 ( .A(n308), .B(n309), .C(n310), .Z(n307) );
  GTECH_XOR2 U157 ( .A(n287), .B(n311), .Z(sum[4]) );
  GTECH_MUX2 U158 ( .A(n312), .B(n313), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U159 ( .A(n314), .B(n315), .Z(n313) );
  GTECH_XNOR2 U160 ( .A(n314), .B(n316), .Z(n312) );
  GTECH_AOI21 U161 ( .A(n317), .B(n318), .C(n319), .Z(n316) );
  GTECH_XOR2 U162 ( .A(a[3]), .B(b[3]), .Z(n314) );
  GTECH_MUX2 U163 ( .A(n320), .B(n321), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U164 ( .A(n322), .B(n323), .Z(n321) );
  GTECH_XOR2 U165 ( .A(n322), .B(n318), .Z(n320) );
  GTECH_OAI21 U166 ( .A(n324), .B(n325), .C(n326), .Z(n318) );
  GTECH_NOT U167 ( .A(n327), .Z(n325) );
  GTECH_AND_NOT U168 ( .A(n317), .B(n319), .Z(n322) );
  GTECH_MUX2 U169 ( .A(n328), .B(n329), .S(n330), .Z(sum[1]) );
  GTECH_AND_NOT U170 ( .A(n326), .B(n324), .Z(n330) );
  GTECH_OAI21 U171 ( .A(cin), .B(n327), .C(n331), .Z(n329) );
  GTECH_NOT U172 ( .A(n332), .Z(n328) );
  GTECH_AOI21 U173 ( .A(n331), .B(cin), .C(n327), .Z(n332) );
  GTECH_MUX2 U174 ( .A(n333), .B(n334), .S(n335), .Z(sum[15]) );
  GTECH_XOR2 U175 ( .A(n336), .B(n337), .Z(n334) );
  GTECH_XNOR2 U176 ( .A(n338), .B(n336), .Z(n333) );
  GTECH_XNOR2 U177 ( .A(a[15]), .B(b[15]), .Z(n336) );
  GTECH_AOI21 U178 ( .A(n339), .B(n340), .C(n341), .Z(n338) );
  GTECH_AOI21 U179 ( .A(n342), .B(a[14]), .C(b[14]), .Z(n341) );
  GTECH_NOT U180 ( .A(n340), .Z(n342) );
  GTECH_NOT U181 ( .A(a[14]), .Z(n339) );
  GTECH_MUX2 U182 ( .A(n343), .B(n344), .S(n335), .Z(sum[14]) );
  GTECH_XOR2 U183 ( .A(n345), .B(n346), .Z(n344) );
  GTECH_XNOR2 U184 ( .A(n345), .B(n340), .Z(n343) );
  GTECH_OA21 U185 ( .A(n347), .B(n348), .C(n349), .Z(n340) );
  GTECH_XOR2 U186 ( .A(a[14]), .B(b[14]), .Z(n345) );
  GTECH_MUX2 U187 ( .A(n350), .B(n351), .S(n335), .Z(sum[13]) );
  GTECH_XNOR2 U188 ( .A(n352), .B(n353), .Z(n351) );
  GTECH_XOR2 U189 ( .A(n354), .B(n352), .Z(n350) );
  GTECH_NOR2 U190 ( .A(n355), .B(n347), .Z(n352) );
  GTECH_OAI21 U191 ( .A(n356), .B(n357), .C(n358), .Z(sum[12]) );
  GTECH_AND2 U192 ( .A(n359), .B(n348), .Z(n356) );
  GTECH_MUX2 U193 ( .A(n360), .B(n361), .S(n284), .Z(sum[11]) );
  GTECH_XOR2 U194 ( .A(n362), .B(n363), .Z(n361) );
  GTECH_XOR2 U195 ( .A(n364), .B(n362), .Z(n360) );
  GTECH_XNOR2 U196 ( .A(n365), .B(b[11]), .Z(n362) );
  GTECH_AOI21 U197 ( .A(n366), .B(n367), .C(n368), .Z(n364) );
  GTECH_AOI21 U198 ( .A(n369), .B(a[10]), .C(b[10]), .Z(n368) );
  GTECH_NOT U199 ( .A(n367), .Z(n369) );
  GTECH_NOT U200 ( .A(a[10]), .Z(n366) );
  GTECH_MUX2 U201 ( .A(n370), .B(n371), .S(n284), .Z(sum[10]) );
  GTECH_NOT U202 ( .A(n277), .Z(n284) );
  GTECH_XNOR2 U203 ( .A(n372), .B(n373), .Z(n371) );
  GTECH_XNOR2 U204 ( .A(n372), .B(n367), .Z(n370) );
  GTECH_AOI21 U205 ( .A(n281), .B(n278), .C(n282), .Z(n367) );
  GTECH_XOR2 U206 ( .A(a[10]), .B(b[10]), .Z(n372) );
  GTECH_XOR2 U207 ( .A(cin), .B(n306), .Z(sum[0]) );
  GTECH_OAI21 U208 ( .A(n374), .B(n357), .C(n358), .Z(cout) );
  GTECH_NAND3 U209 ( .A(n348), .B(n359), .C(n357), .Z(n358) );
  GTECH_NOT U210 ( .A(n354), .Z(n348) );
  GTECH_AND2 U211 ( .A(a[12]), .B(b[12]), .Z(n354) );
  GTECH_NOT U212 ( .A(n335), .Z(n357) );
  GTECH_MUX2 U213 ( .A(n375), .B(n283), .S(n277), .Z(n335) );
  GTECH_MUX2 U214 ( .A(n376), .B(n311), .S(n287), .Z(n277) );
  GTECH_MUX2 U215 ( .A(n377), .B(n378), .S(cin), .Z(n287) );
  GTECH_OA21 U216 ( .A(n308), .B(n309), .C(n310), .Z(n378) );
  GTECH_OAI21 U217 ( .A(a[3]), .B(n315), .C(b[3]), .Z(n310) );
  GTECH_NOT U218 ( .A(n308), .Z(n315) );
  GTECH_NOT U219 ( .A(a[3]), .Z(n309) );
  GTECH_AOI21 U220 ( .A(n317), .B(n323), .C(n319), .Z(n308) );
  GTECH_AND2 U221 ( .A(b[2]), .B(a[2]), .Z(n319) );
  GTECH_OAI21 U222 ( .A(n324), .B(n379), .C(n326), .Z(n323) );
  GTECH_NOT U223 ( .A(n380), .Z(n326) );
  GTECH_AND2 U224 ( .A(b[1]), .B(a[1]), .Z(n380) );
  GTECH_NOR2 U225 ( .A(b[1]), .B(a[1]), .Z(n324) );
  GTECH_OR2 U226 ( .A(a[2]), .B(b[2]), .Z(n317) );
  GTECH_NOT U227 ( .A(n306), .Z(n377) );
  GTECH_NOR2 U228 ( .A(n379), .B(n327), .Z(n306) );
  GTECH_AND2 U229 ( .A(a[0]), .B(b[0]), .Z(n327) );
  GTECH_NOT U230 ( .A(n331), .Z(n379) );
  GTECH_OR2 U231 ( .A(b[0]), .B(a[0]), .Z(n331) );
  GTECH_XNOR2 U232 ( .A(a[4]), .B(b[4]), .Z(n311) );
  GTECH_AOI21 U233 ( .A(n293), .B(a[7]), .C(n381), .Z(n376) );
  GTECH_OA21 U234 ( .A(a[7]), .B(n293), .C(b[7]), .Z(n381) );
  GTECH_OAI21 U235 ( .A(n290), .B(n300), .C(n292), .Z(n293) );
  GTECH_NOT U236 ( .A(n301), .Z(n292) );
  GTECH_AND2 U237 ( .A(b[6]), .B(a[6]), .Z(n301) );
  GTECH_OA21 U238 ( .A(n299), .B(n382), .C(n304), .Z(n300) );
  GTECH_NOT U239 ( .A(n298), .Z(n304) );
  GTECH_AND2 U240 ( .A(a[5]), .B(b[5]), .Z(n298) );
  GTECH_NOR2 U241 ( .A(a[4]), .B(b[4]), .Z(n382) );
  GTECH_NOR2 U242 ( .A(b[5]), .B(a[5]), .Z(n299) );
  GTECH_NOR2 U243 ( .A(b[6]), .B(a[6]), .Z(n290) );
  GTECH_AND_NOT U244 ( .A(n280), .B(n278), .Z(n283) );
  GTECH_AND2 U245 ( .A(a[8]), .B(b[8]), .Z(n278) );
  GTECH_AOI21 U246 ( .A(n365), .B(n383), .C(n384), .Z(n375) );
  GTECH_AOI21 U247 ( .A(n363), .B(a[11]), .C(b[11]), .Z(n384) );
  GTECH_NOT U248 ( .A(n383), .Z(n363) );
  GTECH_AOI21 U249 ( .A(n385), .B(a[10]), .C(n386), .Z(n383) );
  GTECH_OA21 U250 ( .A(a[10]), .B(n385), .C(b[10]), .Z(n386) );
  GTECH_NOT U251 ( .A(n373), .Z(n385) );
  GTECH_AOI21 U252 ( .A(n281), .B(n280), .C(n282), .Z(n373) );
  GTECH_AND2 U253 ( .A(b[9]), .B(a[9]), .Z(n282) );
  GTECH_OR2 U254 ( .A(b[8]), .B(a[8]), .Z(n280) );
  GTECH_OR2 U255 ( .A(a[9]), .B(b[9]), .Z(n281) );
  GTECH_NOT U256 ( .A(a[11]), .Z(n365) );
  GTECH_AOI21 U257 ( .A(n387), .B(a[15]), .C(n388), .Z(n374) );
  GTECH_OA21 U258 ( .A(a[15]), .B(n387), .C(b[15]), .Z(n388) );
  GTECH_NOT U259 ( .A(n337), .Z(n387) );
  GTECH_AOI21 U260 ( .A(n346), .B(a[14]), .C(n389), .Z(n337) );
  GTECH_OA21 U261 ( .A(a[14]), .B(n346), .C(b[14]), .Z(n389) );
  GTECH_OAI21 U262 ( .A(n347), .B(n353), .C(n349), .Z(n346) );
  GTECH_NOT U263 ( .A(n355), .Z(n349) );
  GTECH_AND2 U264 ( .A(b[13]), .B(a[13]), .Z(n355) );
  GTECH_NOT U265 ( .A(n359), .Z(n353) );
  GTECH_OR2 U266 ( .A(b[12]), .B(a[12]), .Z(n359) );
  GTECH_NOR2 U267 ( .A(b[13]), .B(a[13]), .Z(n347) );
endmodule

