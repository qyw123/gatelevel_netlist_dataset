
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n85) );
  GTECH_XNOR2 U78 ( .A(n84), .B(n90), .Z(N154) );
  GTECH_XNOR2 U79 ( .A(n91), .B(n92), .Z(n90) );
  GTECH_NOT U80 ( .A(n86), .Z(n92) );
  GTECH_XNOR2 U81 ( .A(n93), .B(n88), .Z(n86) );
  GTECH_NOT U82 ( .A(n94), .Z(n88) );
  GTECH_NAND2 U83 ( .A(I_b[7]), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U84 ( .A(n89), .Z(n93) );
  GTECH_OAI21 U85 ( .A(n95), .B(n96), .C(n97), .Z(n89) );
  GTECH_OAI21 U86 ( .A(n98), .B(n99), .C(n100), .Z(n97) );
  GTECH_NOT U87 ( .A(n99), .Z(n95) );
  GTECH_NOT U88 ( .A(n87), .Z(n91) );
  GTECH_OAI2N2 U89 ( .A(n101), .B(n102), .C(n103), .D(n104), .Z(n87) );
  GTECH_NAND2 U90 ( .A(n101), .B(n102), .Z(n104) );
  GTECH_NOT U91 ( .A(n105), .Z(n84) );
  GTECH_NAND2 U92 ( .A(n106), .B(n107), .Z(n105) );
  GTECH_NOT U93 ( .A(n108), .Z(n106) );
  GTECH_XNOR2 U94 ( .A(n107), .B(n108), .Z(N153) );
  GTECH_XOR3 U95 ( .A(n109), .B(n101), .C(n103), .Z(n108) );
  GTECH_XOR3 U96 ( .A(n98), .B(n100), .C(n99), .Z(n103) );
  GTECH_OAI21 U97 ( .A(n110), .B(n111), .C(n112), .Z(n99) );
  GTECH_OAI21 U98 ( .A(n113), .B(n114), .C(n115), .Z(n112) );
  GTECH_NOT U99 ( .A(n114), .Z(n110) );
  GTECH_NOT U100 ( .A(n116), .Z(n100) );
  GTECH_NAND2 U101 ( .A(I_b[7]), .B(I_a[6]), .Z(n116) );
  GTECH_NOT U102 ( .A(n96), .Z(n98) );
  GTECH_NAND2 U103 ( .A(I_a[7]), .B(I_b[6]), .Z(n96) );
  GTECH_ADD_ABC U104 ( .A(n117), .B(n118), .C(n119), .COUT(n101) );
  GTECH_NOT U105 ( .A(n120), .Z(n119) );
  GTECH_XNOR2 U106 ( .A(n121), .B(n122), .Z(n118) );
  GTECH_NAND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n122) );
  GTECH_NOT U108 ( .A(n102), .Z(n109) );
  GTECH_NAND2 U109 ( .A(I_a[7]), .B(n123), .Z(n102) );
  GTECH_NOT U110 ( .A(n124), .Z(n107) );
  GTECH_NAND2 U111 ( .A(n125), .B(n126), .Z(n124) );
  GTECH_NOT U112 ( .A(n127), .Z(n126) );
  GTECH_XNOR2 U113 ( .A(n127), .B(n125), .Z(N152) );
  GTECH_XOR4 U114 ( .A(n121), .B(n128), .C(n117), .D(n120), .Z(n125) );
  GTECH_XOR3 U115 ( .A(n113), .B(n115), .C(n114), .Z(n120) );
  GTECH_OAI21 U116 ( .A(n129), .B(n130), .C(n131), .Z(n114) );
  GTECH_OAI21 U117 ( .A(n132), .B(n133), .C(n134), .Z(n131) );
  GTECH_NOT U118 ( .A(n133), .Z(n129) );
  GTECH_NOT U119 ( .A(n135), .Z(n115) );
  GTECH_NAND2 U120 ( .A(I_b[7]), .B(I_a[5]), .Z(n135) );
  GTECH_NOT U121 ( .A(n111), .Z(n113) );
  GTECH_NAND2 U122 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_ADD_ABC U123 ( .A(n136), .B(n137), .C(n138), .COUT(n117) );
  GTECH_NOT U124 ( .A(n139), .Z(n138) );
  GTECH_XOR3 U125 ( .A(n140), .B(n141), .C(n142), .Z(n137) );
  GTECH_AND2 U126 ( .A(I_a[7]), .B(I_b[5]), .Z(n128) );
  GTECH_NOT U127 ( .A(n123), .Z(n121) );
  GTECH_OAI21 U128 ( .A(n142), .B(n143), .C(n144), .Z(n123) );
  GTECH_OAI21 U129 ( .A(n140), .B(n145), .C(n141), .Z(n144) );
  GTECH_NOT U130 ( .A(n143), .Z(n140) );
  GTECH_NOT U131 ( .A(n145), .Z(n142) );
  GTECH_ADD_ABC U132 ( .A(n146), .B(n147), .C(n148), .COUT(n127) );
  GTECH_NOT U133 ( .A(n149), .Z(n148) );
  GTECH_OA22 U134 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n147) );
  GTECH_OA21 U135 ( .A(n154), .B(n155), .C(n156), .Z(n146) );
  GTECH_XOR3 U136 ( .A(n157), .B(n149), .C(n158), .Z(N151) );
  GTECH_OA21 U137 ( .A(n154), .B(n155), .C(n156), .Z(n158) );
  GTECH_OAI21 U138 ( .A(n159), .B(n160), .C(n161), .Z(n156) );
  GTECH_XOR3 U139 ( .A(n139), .B(n136), .C(n162), .Z(n149) );
  GTECH_XOR3 U140 ( .A(n141), .B(n145), .C(n143), .Z(n162) );
  GTECH_NAND2 U141 ( .A(I_a[7]), .B(I_b[4]), .Z(n143) );
  GTECH_OAI21 U142 ( .A(n163), .B(n164), .C(n165), .Z(n145) );
  GTECH_OAI21 U143 ( .A(n166), .B(n167), .C(n168), .Z(n165) );
  GTECH_NOT U144 ( .A(n169), .Z(n141) );
  GTECH_NAND2 U145 ( .A(I_a[6]), .B(I_b[5]), .Z(n169) );
  GTECH_ADD_ABC U146 ( .A(n170), .B(n171), .C(n172), .COUT(n136) );
  GTECH_NOT U147 ( .A(n173), .Z(n172) );
  GTECH_XOR3 U148 ( .A(n166), .B(n168), .C(n163), .Z(n171) );
  GTECH_NOT U149 ( .A(n167), .Z(n163) );
  GTECH_NOT U150 ( .A(n164), .Z(n166) );
  GTECH_XOR3 U151 ( .A(n132), .B(n134), .C(n133), .Z(n139) );
  GTECH_OAI21 U152 ( .A(n174), .B(n175), .C(n176), .Z(n133) );
  GTECH_OAI21 U153 ( .A(n177), .B(n178), .C(n179), .Z(n176) );
  GTECH_NOT U154 ( .A(n178), .Z(n174) );
  GTECH_NOT U155 ( .A(n180), .Z(n134) );
  GTECH_NAND2 U156 ( .A(I_b[7]), .B(I_a[4]), .Z(n180) );
  GTECH_NOT U157 ( .A(n130), .Z(n132) );
  GTECH_NAND2 U158 ( .A(I_b[6]), .B(I_a[5]), .Z(n130) );
  GTECH_OA22 U159 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n157) );
  GTECH_NOT U160 ( .A(I_a[7]), .Z(n151) );
  GTECH_XOR3 U161 ( .A(n154), .B(n159), .C(n181), .Z(N150) );
  GTECH_NOT U162 ( .A(n161), .Z(n181) );
  GTECH_XOR3 U163 ( .A(n173), .B(n170), .C(n182), .Z(n161) );
  GTECH_XOR3 U164 ( .A(n168), .B(n167), .C(n164), .Z(n182) );
  GTECH_NAND2 U165 ( .A(I_a[6]), .B(I_b[4]), .Z(n164) );
  GTECH_OAI21 U166 ( .A(n183), .B(n184), .C(n185), .Z(n167) );
  GTECH_OAI21 U167 ( .A(n186), .B(n187), .C(n188), .Z(n185) );
  GTECH_NOT U168 ( .A(n189), .Z(n168) );
  GTECH_NAND2 U169 ( .A(I_a[5]), .B(I_b[5]), .Z(n189) );
  GTECH_ADD_ABC U170 ( .A(n190), .B(n191), .C(n192), .COUT(n170) );
  GTECH_NOT U171 ( .A(n193), .Z(n192) );
  GTECH_XOR3 U172 ( .A(n186), .B(n188), .C(n183), .Z(n191) );
  GTECH_NOT U173 ( .A(n187), .Z(n183) );
  GTECH_NOT U174 ( .A(n184), .Z(n186) );
  GTECH_XOR3 U175 ( .A(n177), .B(n179), .C(n178), .Z(n173) );
  GTECH_OAI21 U176 ( .A(n194), .B(n195), .C(n196), .Z(n178) );
  GTECH_OAI21 U177 ( .A(n197), .B(n198), .C(n199), .Z(n196) );
  GTECH_NOT U178 ( .A(n198), .Z(n194) );
  GTECH_NOT U179 ( .A(n200), .Z(n179) );
  GTECH_NAND2 U180 ( .A(I_b[7]), .B(I_a[3]), .Z(n200) );
  GTECH_NOT U181 ( .A(n175), .Z(n177) );
  GTECH_NAND2 U182 ( .A(I_b[6]), .B(I_a[4]), .Z(n175) );
  GTECH_NOT U183 ( .A(n155), .Z(n159) );
  GTECH_XNOR2 U184 ( .A(n152), .B(n153), .Z(n155) );
  GTECH_XNOR2 U185 ( .A(n150), .B(n201), .Z(n153) );
  GTECH_NAND2 U186 ( .A(I_a[7]), .B(I_b[3]), .Z(n201) );
  GTECH_OA21 U187 ( .A(n202), .B(n203), .C(n204), .Z(n150) );
  GTECH_OAI21 U188 ( .A(n205), .B(n206), .C(n207), .Z(n204) );
  GTECH_NOT U189 ( .A(n206), .Z(n203) );
  GTECH_AOI2N2 U190 ( .A(n208), .B(n209), .C(n210), .D(n211), .Z(n152) );
  GTECH_NAND2 U191 ( .A(n210), .B(n211), .Z(n209) );
  GTECH_NOT U192 ( .A(n160), .Z(n154) );
  GTECH_OAI2N2 U193 ( .A(n212), .B(n213), .C(n214), .D(n215), .Z(n160) );
  GTECH_NAND2 U194 ( .A(n212), .B(n213), .Z(n215) );
  GTECH_XOR3 U195 ( .A(n212), .B(n216), .C(n217), .Z(N149) );
  GTECH_NOT U196 ( .A(n214), .Z(n217) );
  GTECH_XOR3 U197 ( .A(n193), .B(n190), .C(n218), .Z(n214) );
  GTECH_XOR3 U198 ( .A(n188), .B(n187), .C(n184), .Z(n218) );
  GTECH_NAND2 U199 ( .A(I_a[5]), .B(I_b[4]), .Z(n184) );
  GTECH_OAI21 U200 ( .A(n219), .B(n220), .C(n221), .Z(n187) );
  GTECH_OAI21 U201 ( .A(n222), .B(n223), .C(n224), .Z(n221) );
  GTECH_NOT U202 ( .A(n225), .Z(n188) );
  GTECH_NAND2 U203 ( .A(I_b[5]), .B(I_a[4]), .Z(n225) );
  GTECH_ADD_ABC U204 ( .A(n226), .B(n227), .C(n228), .COUT(n190) );
  GTECH_XOR3 U205 ( .A(n222), .B(n224), .C(n219), .Z(n227) );
  GTECH_NOT U206 ( .A(n223), .Z(n219) );
  GTECH_OA21 U207 ( .A(n229), .B(n230), .C(n231), .Z(n226) );
  GTECH_XOR3 U208 ( .A(n197), .B(n199), .C(n198), .Z(n193) );
  GTECH_OAI21 U209 ( .A(n232), .B(n233), .C(n234), .Z(n198) );
  GTECH_NOT U210 ( .A(n235), .Z(n199) );
  GTECH_NAND2 U211 ( .A(I_b[7]), .B(I_a[2]), .Z(n235) );
  GTECH_NOT U212 ( .A(n195), .Z(n197) );
  GTECH_NAND2 U213 ( .A(I_b[6]), .B(I_a[3]), .Z(n195) );
  GTECH_NOT U214 ( .A(n213), .Z(n216) );
  GTECH_XOR3 U215 ( .A(n236), .B(n210), .C(n208), .Z(n213) );
  GTECH_XOR3 U216 ( .A(n205), .B(n207), .C(n206), .Z(n208) );
  GTECH_OAI21 U217 ( .A(n237), .B(n238), .C(n239), .Z(n206) );
  GTECH_OAI21 U218 ( .A(n240), .B(n241), .C(n242), .Z(n239) );
  GTECH_NOT U219 ( .A(n241), .Z(n237) );
  GTECH_NOT U220 ( .A(n243), .Z(n207) );
  GTECH_NAND2 U221 ( .A(I_a[6]), .B(I_b[3]), .Z(n243) );
  GTECH_NOT U222 ( .A(n202), .Z(n205) );
  GTECH_NAND2 U223 ( .A(I_a[7]), .B(I_b[2]), .Z(n202) );
  GTECH_ADD_ABC U224 ( .A(n244), .B(n245), .C(n246), .COUT(n210) );
  GTECH_XNOR2 U225 ( .A(n247), .B(n248), .Z(n245) );
  GTECH_NAND2 U226 ( .A(I_a[7]), .B(I_b[1]), .Z(n248) );
  GTECH_NOT U227 ( .A(n211), .Z(n236) );
  GTECH_NAND2 U228 ( .A(I_a[7]), .B(n249), .Z(n211) );
  GTECH_ADD_ABC U229 ( .A(n250), .B(n251), .C(n252), .COUT(n212) );
  GTECH_XOR3 U230 ( .A(n244), .B(n253), .C(n246), .Z(n251) );
  GTECH_NOT U231 ( .A(n254), .Z(n246) );
  GTECH_XOR3 U232 ( .A(n255), .B(n252), .C(n250), .Z(N148) );
  GTECH_ADD_ABC U233 ( .A(n256), .B(n257), .C(n258), .COUT(n250) );
  GTECH_NOT U234 ( .A(n259), .Z(n258) );
  GTECH_XOR3 U235 ( .A(n260), .B(n261), .C(n262), .Z(n257) );
  GTECH_NOT U236 ( .A(n263), .Z(n261) );
  GTECH_XOR3 U237 ( .A(n264), .B(n228), .C(n265), .Z(n252) );
  GTECH_OAI21 U238 ( .A(n229), .B(n230), .C(n231), .Z(n265) );
  GTECH_OAI21 U239 ( .A(n266), .B(n267), .C(n268), .Z(n231) );
  GTECH_NOT U240 ( .A(n229), .Z(n267) );
  GTECH_XOR3 U241 ( .A(n269), .B(n270), .C(n234), .Z(n228) );
  GTECH_NAND3 U242 ( .A(I_b[7]), .B(I_a[0]), .C(n271), .Z(n234) );
  GTECH_NOT U243 ( .A(n233), .Z(n270) );
  GTECH_NAND2 U244 ( .A(I_b[7]), .B(I_a[1]), .Z(n233) );
  GTECH_NOT U245 ( .A(n232), .Z(n269) );
  GTECH_NAND2 U246 ( .A(I_b[6]), .B(I_a[2]), .Z(n232) );
  GTECH_XOR3 U247 ( .A(n224), .B(n223), .C(n222), .Z(n264) );
  GTECH_NOT U248 ( .A(n220), .Z(n222) );
  GTECH_NAND2 U249 ( .A(I_b[4]), .B(I_a[4]), .Z(n220) );
  GTECH_OAI21 U250 ( .A(n272), .B(n273), .C(n274), .Z(n223) );
  GTECH_OAI21 U251 ( .A(n275), .B(n276), .C(n277), .Z(n274) );
  GTECH_NOT U252 ( .A(n276), .Z(n272) );
  GTECH_NOT U253 ( .A(n278), .Z(n224) );
  GTECH_NAND2 U254 ( .A(I_b[5]), .B(I_a[3]), .Z(n278) );
  GTECH_XOR3 U255 ( .A(n253), .B(n254), .C(n244), .Z(n255) );
  GTECH_ADD_ABC U256 ( .A(n260), .B(n279), .C(n262), .COUT(n244) );
  GTECH_NOT U257 ( .A(n280), .Z(n262) );
  GTECH_XOR3 U258 ( .A(n281), .B(n282), .C(n283), .Z(n279) );
  GTECH_XOR3 U259 ( .A(n240), .B(n242), .C(n241), .Z(n254) );
  GTECH_OAI21 U260 ( .A(n284), .B(n285), .C(n286), .Z(n241) );
  GTECH_OAI21 U261 ( .A(n287), .B(n288), .C(n289), .Z(n286) );
  GTECH_NOT U262 ( .A(n288), .Z(n284) );
  GTECH_NOT U263 ( .A(n290), .Z(n242) );
  GTECH_NAND2 U264 ( .A(I_a[5]), .B(I_b[3]), .Z(n290) );
  GTECH_NOT U265 ( .A(n238), .Z(n240) );
  GTECH_NAND2 U266 ( .A(I_a[6]), .B(I_b[2]), .Z(n238) );
  GTECH_XNOR2 U267 ( .A(n247), .B(n291), .Z(n253) );
  GTECH_NAND2 U268 ( .A(I_a[7]), .B(I_b[1]), .Z(n291) );
  GTECH_NOT U269 ( .A(n249), .Z(n247) );
  GTECH_OAI21 U270 ( .A(n283), .B(n292), .C(n293), .Z(n249) );
  GTECH_OAI21 U271 ( .A(n281), .B(n294), .C(n282), .Z(n293) );
  GTECH_NOT U272 ( .A(n294), .Z(n283) );
  GTECH_XOR3 U273 ( .A(n259), .B(n256), .C(n295), .Z(N147) );
  GTECH_XOR3 U274 ( .A(n280), .B(n260), .C(n263), .Z(n295) );
  GTECH_XOR3 U275 ( .A(n281), .B(n282), .C(n294), .Z(n263) );
  GTECH_OAI21 U276 ( .A(n296), .B(n297), .C(n298), .Z(n294) );
  GTECH_OAI21 U277 ( .A(n299), .B(n300), .C(n301), .Z(n298) );
  GTECH_NOT U278 ( .A(n302), .Z(n282) );
  GTECH_NAND2 U279 ( .A(I_a[6]), .B(I_b[1]), .Z(n302) );
  GTECH_NOT U280 ( .A(n292), .Z(n281) );
  GTECH_NAND2 U281 ( .A(I_a[7]), .B(I_b[0]), .Z(n292) );
  GTECH_ADD_ABC U282 ( .A(n303), .B(n304), .C(n305), .COUT(n260) );
  GTECH_XOR3 U283 ( .A(n299), .B(n301), .C(n296), .Z(n304) );
  GTECH_NOT U284 ( .A(n300), .Z(n296) );
  GTECH_XOR3 U285 ( .A(n287), .B(n289), .C(n288), .Z(n280) );
  GTECH_OAI21 U286 ( .A(n306), .B(n307), .C(n308), .Z(n288) );
  GTECH_OAI21 U287 ( .A(n309), .B(n310), .C(n311), .Z(n308) );
  GTECH_NOT U288 ( .A(n310), .Z(n306) );
  GTECH_NOT U289 ( .A(n312), .Z(n289) );
  GTECH_NAND2 U290 ( .A(I_b[3]), .B(I_a[4]), .Z(n312) );
  GTECH_NOT U291 ( .A(n285), .Z(n287) );
  GTECH_NAND2 U292 ( .A(I_a[5]), .B(I_b[2]), .Z(n285) );
  GTECH_ADD_ABC U293 ( .A(n313), .B(n314), .C(n315), .COUT(n256) );
  GTECH_XOR3 U294 ( .A(n303), .B(n316), .C(n305), .Z(n314) );
  GTECH_NOT U295 ( .A(n317), .Z(n305) );
  GTECH_OA21 U296 ( .A(n318), .B(n319), .C(n320), .Z(n313) );
  GTECH_XOR3 U297 ( .A(n268), .B(n230), .C(n229), .Z(n259) );
  GTECH_XNOR2 U298 ( .A(n271), .B(n321), .Z(n229) );
  GTECH_AND2 U299 ( .A(I_b[7]), .B(I_a[0]), .Z(n321) );
  GTECH_NOT U300 ( .A(n322), .Z(n271) );
  GTECH_NAND2 U301 ( .A(I_b[6]), .B(I_a[1]), .Z(n322) );
  GTECH_NOT U302 ( .A(n266), .Z(n230) );
  GTECH_XOR3 U303 ( .A(n275), .B(n277), .C(n276), .Z(n266) );
  GTECH_OAI21 U304 ( .A(n323), .B(n324), .C(n325), .Z(n276) );
  GTECH_NOT U305 ( .A(n326), .Z(n277) );
  GTECH_NAND2 U306 ( .A(I_b[5]), .B(I_a[2]), .Z(n326) );
  GTECH_NOT U307 ( .A(n273), .Z(n275) );
  GTECH_NAND2 U308 ( .A(I_b[4]), .B(I_a[3]), .Z(n273) );
  GTECH_NOT U309 ( .A(n327), .Z(n268) );
  GTECH_NAND3 U310 ( .A(I_a[0]), .B(n328), .C(I_b[6]), .Z(n327) );
  GTECH_XOR3 U311 ( .A(n329), .B(n315), .C(n330), .Z(N146) );
  GTECH_OA21 U312 ( .A(n318), .B(n319), .C(n320), .Z(n330) );
  GTECH_OAI21 U313 ( .A(n331), .B(n332), .C(n333), .Z(n320) );
  GTECH_NOT U314 ( .A(n318), .Z(n332) );
  GTECH_XNOR2 U315 ( .A(n334), .B(n328), .Z(n315) );
  GTECH_NOT U316 ( .A(n335), .Z(n328) );
  GTECH_XOR3 U317 ( .A(n336), .B(n337), .C(n325), .Z(n335) );
  GTECH_NAND3 U318 ( .A(I_b[5]), .B(I_a[0]), .C(n338), .Z(n325) );
  GTECH_NOT U319 ( .A(n324), .Z(n337) );
  GTECH_NAND2 U320 ( .A(I_b[5]), .B(I_a[1]), .Z(n324) );
  GTECH_NOT U321 ( .A(n323), .Z(n336) );
  GTECH_NAND2 U322 ( .A(I_b[4]), .B(I_a[2]), .Z(n323) );
  GTECH_AND2 U323 ( .A(I_b[6]), .B(I_a[0]), .Z(n334) );
  GTECH_XOR3 U324 ( .A(n316), .B(n317), .C(n303), .Z(n329) );
  GTECH_ADD_ABC U325 ( .A(n339), .B(n340), .C(n341), .COUT(n303) );
  GTECH_NOT U326 ( .A(n342), .Z(n341) );
  GTECH_XOR3 U327 ( .A(n343), .B(n344), .C(n345), .Z(n340) );
  GTECH_XOR3 U328 ( .A(n309), .B(n311), .C(n310), .Z(n317) );
  GTECH_OAI21 U329 ( .A(n346), .B(n347), .C(n348), .Z(n310) );
  GTECH_OAI21 U330 ( .A(n349), .B(n350), .C(n351), .Z(n348) );
  GTECH_NOT U331 ( .A(n350), .Z(n346) );
  GTECH_NOT U332 ( .A(n352), .Z(n311) );
  GTECH_NAND2 U333 ( .A(I_b[3]), .B(I_a[3]), .Z(n352) );
  GTECH_NOT U334 ( .A(n307), .Z(n309) );
  GTECH_NAND2 U335 ( .A(I_b[2]), .B(I_a[4]), .Z(n307) );
  GTECH_NOT U336 ( .A(n353), .Z(n316) );
  GTECH_XOR3 U337 ( .A(n299), .B(n301), .C(n300), .Z(n353) );
  GTECH_OAI21 U338 ( .A(n345), .B(n354), .C(n355), .Z(n300) );
  GTECH_OAI21 U339 ( .A(n343), .B(n356), .C(n344), .Z(n355) );
  GTECH_NOT U340 ( .A(n354), .Z(n343) );
  GTECH_NOT U341 ( .A(n356), .Z(n345) );
  GTECH_NOT U342 ( .A(n357), .Z(n301) );
  GTECH_NAND2 U343 ( .A(I_a[5]), .B(I_b[1]), .Z(n357) );
  GTECH_NOT U344 ( .A(n297), .Z(n299) );
  GTECH_NAND2 U345 ( .A(I_a[6]), .B(I_b[0]), .Z(n297) );
  GTECH_XOR3 U346 ( .A(n333), .B(n319), .C(n318), .Z(N145) );
  GTECH_XNOR2 U347 ( .A(n338), .B(n358), .Z(n318) );
  GTECH_AND2 U348 ( .A(I_b[5]), .B(I_a[0]), .Z(n358) );
  GTECH_NOT U349 ( .A(n359), .Z(n338) );
  GTECH_NAND2 U350 ( .A(I_b[4]), .B(I_a[1]), .Z(n359) );
  GTECH_NOT U351 ( .A(n331), .Z(n319) );
  GTECH_XOR3 U352 ( .A(n342), .B(n339), .C(n360), .Z(n331) );
  GTECH_XOR3 U353 ( .A(n344), .B(n356), .C(n354), .Z(n360) );
  GTECH_NAND2 U354 ( .A(I_a[5]), .B(I_b[0]), .Z(n354) );
  GTECH_OAI21 U355 ( .A(n361), .B(n362), .C(n363), .Z(n356) );
  GTECH_OAI21 U356 ( .A(n364), .B(n365), .C(n366), .Z(n363) );
  GTECH_NOT U357 ( .A(n367), .Z(n344) );
  GTECH_NAND2 U358 ( .A(I_a[4]), .B(I_b[1]), .Z(n367) );
  GTECH_ADD_ABC U359 ( .A(n368), .B(n369), .C(n370), .COUT(n339) );
  GTECH_XOR3 U360 ( .A(n364), .B(n366), .C(n361), .Z(n369) );
  GTECH_NOT U361 ( .A(n365), .Z(n361) );
  GTECH_OA21 U362 ( .A(n371), .B(n372), .C(n373), .Z(n368) );
  GTECH_XOR3 U363 ( .A(n349), .B(n351), .C(n350), .Z(n342) );
  GTECH_OAI21 U364 ( .A(n374), .B(n375), .C(n376), .Z(n350) );
  GTECH_NOT U365 ( .A(n377), .Z(n351) );
  GTECH_NAND2 U366 ( .A(I_b[3]), .B(I_a[2]), .Z(n377) );
  GTECH_NOT U367 ( .A(n347), .Z(n349) );
  GTECH_NAND2 U368 ( .A(I_b[2]), .B(I_a[3]), .Z(n347) );
  GTECH_NOT U369 ( .A(n378), .Z(n333) );
  GTECH_NAND3 U370 ( .A(I_a[0]), .B(n379), .C(I_b[4]), .Z(n378) );
  GTECH_NOT U371 ( .A(n380), .Z(n379) );
  GTECH_XNOR2 U372 ( .A(n381), .B(n380), .Z(N144) );
  GTECH_XOR3 U373 ( .A(n382), .B(n370), .C(n383), .Z(n380) );
  GTECH_OAI21 U374 ( .A(n371), .B(n372), .C(n373), .Z(n383) );
  GTECH_OAI21 U375 ( .A(n384), .B(n385), .C(n386), .Z(n373) );
  GTECH_NOT U376 ( .A(n371), .Z(n385) );
  GTECH_XOR3 U377 ( .A(n387), .B(n388), .C(n376), .Z(n370) );
  GTECH_NAND3 U378 ( .A(I_b[3]), .B(I_a[0]), .C(n389), .Z(n376) );
  GTECH_NOT U379 ( .A(n375), .Z(n388) );
  GTECH_NAND2 U380 ( .A(I_b[3]), .B(I_a[1]), .Z(n375) );
  GTECH_NOT U381 ( .A(n374), .Z(n387) );
  GTECH_NAND2 U382 ( .A(I_b[2]), .B(I_a[2]), .Z(n374) );
  GTECH_XOR3 U383 ( .A(n366), .B(n365), .C(n364), .Z(n382) );
  GTECH_NOT U384 ( .A(n362), .Z(n364) );
  GTECH_NAND2 U385 ( .A(I_a[4]), .B(I_b[0]), .Z(n362) );
  GTECH_OAI21 U386 ( .A(n390), .B(n391), .C(n392), .Z(n365) );
  GTECH_OAI21 U387 ( .A(n393), .B(n394), .C(n395), .Z(n392) );
  GTECH_NOT U388 ( .A(n394), .Z(n390) );
  GTECH_NOT U389 ( .A(n396), .Z(n366) );
  GTECH_NAND2 U390 ( .A(I_a[3]), .B(I_b[1]), .Z(n396) );
  GTECH_AND2 U391 ( .A(I_b[4]), .B(I_a[0]), .Z(n381) );
  GTECH_XOR3 U392 ( .A(n386), .B(n372), .C(n371), .Z(N143) );
  GTECH_XNOR2 U393 ( .A(n389), .B(n397), .Z(n371) );
  GTECH_AND2 U394 ( .A(I_b[3]), .B(I_a[0]), .Z(n397) );
  GTECH_NOT U395 ( .A(n398), .Z(n389) );
  GTECH_NAND2 U396 ( .A(I_b[2]), .B(I_a[1]), .Z(n398) );
  GTECH_NOT U397 ( .A(n384), .Z(n372) );
  GTECH_XOR3 U398 ( .A(n393), .B(n395), .C(n394), .Z(n384) );
  GTECH_OAI21 U399 ( .A(n399), .B(n400), .C(n401), .Z(n394) );
  GTECH_NOT U400 ( .A(n402), .Z(n395) );
  GTECH_NAND2 U401 ( .A(I_b[1]), .B(I_a[2]), .Z(n402) );
  GTECH_NOT U402 ( .A(n391), .Z(n393) );
  GTECH_NAND2 U403 ( .A(I_b[0]), .B(I_a[3]), .Z(n391) );
  GTECH_NOT U404 ( .A(n403), .Z(n386) );
  GTECH_NAND3 U405 ( .A(I_a[0]), .B(n404), .C(I_b[2]), .Z(n403) );
  GTECH_NOT U406 ( .A(n405), .Z(n404) );
  GTECH_XNOR2 U407 ( .A(n406), .B(n405), .Z(N142) );
  GTECH_XOR3 U408 ( .A(n407), .B(n408), .C(n401), .Z(n405) );
  GTECH_NAND3 U409 ( .A(n409), .B(I_b[1]), .C(I_a[0]), .Z(n401) );
  GTECH_NOT U410 ( .A(n399), .Z(n408) );
  GTECH_NAND2 U411 ( .A(I_a[1]), .B(I_b[1]), .Z(n399) );
  GTECH_NOT U412 ( .A(n400), .Z(n407) );
  GTECH_NAND2 U413 ( .A(I_b[0]), .B(I_a[2]), .Z(n400) );
  GTECH_AND2 U414 ( .A(I_b[2]), .B(I_a[0]), .Z(n406) );
  GTECH_XNOR2 U415 ( .A(n409), .B(n410), .Z(N141) );
  GTECH_NAND2 U416 ( .A(I_a[0]), .B(I_b[1]), .Z(n410) );
  GTECH_NOT U417 ( .A(n411), .Z(n409) );
  GTECH_NAND2 U418 ( .A(I_a[1]), .B(I_b[0]), .Z(n411) );
  GTECH_AND2 U419 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

