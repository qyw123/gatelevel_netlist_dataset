
module carry_select_adder8 ( a, b, cin, cout, sum );
  input [7:0] a;
  input [7:0] b;
  output [7:0] sum;
  input cin;
  output cout;
  wire   n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187;

  GTECH_MUX2 U66 ( .A(n135), .B(n136), .S(n137), .Z(sum[7]) );
  GTECH_XOR2 U67 ( .A(n138), .B(n139), .Z(n136) );
  GTECH_OA21 U68 ( .A(n140), .B(n141), .C(n142), .Z(n139) );
  GTECH_XOR2 U69 ( .A(n138), .B(n143), .Z(n135) );
  GTECH_XNOR2 U70 ( .A(n144), .B(n145), .Z(n138) );
  GTECH_MUX2 U71 ( .A(n146), .B(n147), .S(n137), .Z(sum[6]) );
  GTECH_XNOR2 U72 ( .A(n141), .B(n148), .Z(n147) );
  GTECH_OA21 U73 ( .A(n149), .B(n150), .C(n151), .Z(n141) );
  GTECH_XNOR2 U74 ( .A(n148), .B(n152), .Z(n146) );
  GTECH_AND_NOT U75 ( .A(n142), .B(n140), .Z(n148) );
  GTECH_MUX2 U76 ( .A(n153), .B(n154), .S(n155), .Z(sum[5]) );
  GTECH_AOI21 U77 ( .A(n149), .B(n137), .C(n156), .Z(n155) );
  GTECH_OR_NOT U78 ( .A(n150), .B(n151), .Z(n154) );
  GTECH_XOR2 U79 ( .A(b[5]), .B(a[5]), .Z(n153) );
  GTECH_OR_NOT U80 ( .A(n157), .B(n158), .Z(sum[4]) );
  GTECH_AO21 U81 ( .A(n149), .B(n159), .C(n137), .Z(n158) );
  GTECH_MUX2 U82 ( .A(n160), .B(n161), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U83 ( .A(n162), .B(n163), .Z(n161) );
  GTECH_XOR2 U84 ( .A(n162), .B(n164), .Z(n160) );
  GTECH_AOI21 U85 ( .A(n165), .B(n166), .C(n167), .Z(n164) );
  GTECH_XNOR2 U86 ( .A(a[3]), .B(b[3]), .Z(n162) );
  GTECH_MUX2 U87 ( .A(n168), .B(n169), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U88 ( .A(n170), .B(n171), .Z(n169) );
  GTECH_XOR2 U89 ( .A(n166), .B(n171), .Z(n168) );
  GTECH_AND_NOT U90 ( .A(n165), .B(n167), .Z(n171) );
  GTECH_OR_NOT U91 ( .A(n172), .B(n173), .Z(n166) );
  GTECH_NAND3 U92 ( .A(b[0]), .B(n174), .C(a[0]), .Z(n173) );
  GTECH_MUX2 U93 ( .A(n175), .B(n176), .S(cin), .Z(sum[1]) );
  GTECH_XOR2 U94 ( .A(n177), .B(n178), .Z(n176) );
  GTECH_XOR2 U95 ( .A(n177), .B(n179), .Z(n175) );
  GTECH_AND2 U96 ( .A(a[0]), .B(b[0]), .Z(n179) );
  GTECH_AND_NOT U97 ( .A(n174), .B(n172), .Z(n177) );
  GTECH_XNOR2 U98 ( .A(cin), .B(n180), .Z(sum[0]) );
  GTECH_AO21 U99 ( .A(n181), .B(n182), .C(n157), .Z(cout) );
  GTECH_AND3 U100 ( .A(n159), .B(n149), .C(n137), .Z(n157) );
  GTECH_NAND2 U101 ( .A(b[4]), .B(a[4]), .Z(n149) );
  GTECH_OAI22 U102 ( .A(n143), .B(n144), .C(n183), .D(n145), .Z(n182) );
  GTECH_NOT U103 ( .A(b[7]), .Z(n145) );
  GTECH_AND_NOT U104 ( .A(n143), .B(a[7]), .Z(n183) );
  GTECH_NOT U105 ( .A(a[7]), .Z(n144) );
  GTECH_OA21 U106 ( .A(n140), .B(n152), .C(n142), .Z(n143) );
  GTECH_OR_NOT U107 ( .A(n184), .B(b[6]), .Z(n142) );
  GTECH_OA21 U108 ( .A(n156), .B(n150), .C(n151), .Z(n152) );
  GTECH_NAND2 U109 ( .A(b[5]), .B(a[5]), .Z(n151) );
  GTECH_NOT U110 ( .A(n185), .Z(n150) );
  GTECH_OR2 U111 ( .A(a[5]), .B(b[5]), .Z(n185) );
  GTECH_NOT U112 ( .A(n159), .Z(n156) );
  GTECH_OR2 U113 ( .A(a[4]), .B(b[4]), .Z(n159) );
  GTECH_AND_NOT U114 ( .A(n184), .B(b[6]), .Z(n140) );
  GTECH_NOT U115 ( .A(a[6]), .Z(n184) );
  GTECH_NOT U116 ( .A(n137), .Z(n181) );
  GTECH_MUX2 U117 ( .A(n180), .B(n186), .S(cin), .Z(n137) );
  GTECH_AOI21 U118 ( .A(n163), .B(a[3]), .C(n187), .Z(n186) );
  GTECH_OA21 U119 ( .A(n163), .B(a[3]), .C(b[3]), .Z(n187) );
  GTECH_AO21 U120 ( .A(n165), .B(n170), .C(n167), .Z(n163) );
  GTECH_AND2 U121 ( .A(b[2]), .B(a[2]), .Z(n167) );
  GTECH_AO21 U122 ( .A(n174), .B(n178), .C(n172), .Z(n170) );
  GTECH_AND2 U123 ( .A(b[1]), .B(a[1]), .Z(n172) );
  GTECH_OR2 U124 ( .A(a[0]), .B(b[0]), .Z(n178) );
  GTECH_OR2 U125 ( .A(a[1]), .B(b[1]), .Z(n174) );
  GTECH_OR2 U126 ( .A(b[2]), .B(a[2]), .Z(n165) );
  GTECH_XNOR2 U127 ( .A(a[0]), .B(b[0]), .Z(n180) );
endmodule

