
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_XOR2 U75 ( .A(n83), .B(n84), .Z(N155) );
  GTECH_AND2 U76 ( .A(n85), .B(n86), .Z(n84) );
  GTECH_OAI22 U77 ( .A(n87), .B(n88), .C(n89), .D(n90), .Z(n83) );
  GTECH_XOR2 U78 ( .A(n85), .B(n86), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n86) );
  GTECH_XOR2 U80 ( .A(n89), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n90), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n90) );
  GTECH_OR_NOT U83 ( .A(n97), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n88), .B(n98), .Z(n89) );
  GTECH_NOT U85 ( .A(n87), .Z(n98) );
  GTECH_OAI22 U86 ( .A(n99), .B(n100), .C(n101), .D(n102), .Z(n87) );
  GTECH_NOR2 U87 ( .A(n103), .B(n104), .Z(n99) );
  GTECH_OR_NOT U88 ( .A(n105), .B(I_b[7]), .Z(n88) );
  GTECH_NOT U89 ( .A(n106), .Z(n85) );
  GTECH_OR_NOT U90 ( .A(n107), .B(n108), .Z(n106) );
  GTECH_XOR2 U91 ( .A(n109), .B(n108), .Z(N153) );
  GTECH_NOT U92 ( .A(n110), .Z(n108) );
  GTECH_XOR3 U93 ( .A(n93), .B(n95), .C(n94), .Z(n110) );
  GTECH_XOR3 U94 ( .A(n101), .B(n102), .C(n100), .Z(n94) );
  GTECH_OAI21 U95 ( .A(n111), .B(n112), .C(n113), .Z(n100) );
  GTECH_OAI21 U96 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_NOT U97 ( .A(n104), .Z(n102) );
  GTECH_OR_NOT U98 ( .A(n117), .B(I_a[7]), .Z(n104) );
  GTECH_NOT U99 ( .A(I_b[6]), .Z(n117) );
  GTECH_NOT U100 ( .A(n103), .Z(n101) );
  GTECH_OR_NOT U101 ( .A(n118), .B(I_b[7]), .Z(n103) );
  GTECH_AOI2N2 U102 ( .A(n119), .B(n120), .C(n121), .D(n122), .Z(n95) );
  GTECH_OR_NOT U103 ( .A(n123), .B(n121), .Z(n120) );
  GTECH_NOT U104 ( .A(n97), .Z(n93) );
  GTECH_OR_NOT U105 ( .A(n105), .B(n124), .Z(n97) );
  GTECH_NOT U106 ( .A(n107), .Z(n109) );
  GTECH_OR_NOT U107 ( .A(n125), .B(n126), .Z(n107) );
  GTECH_NOT U108 ( .A(n127), .Z(n126) );
  GTECH_XOR2 U109 ( .A(n127), .B(n125), .Z(N152) );
  GTECH_AOI22 U110 ( .A(n128), .B(n129), .C(n130), .D(n131), .Z(n125) );
  GTECH_OR2 U111 ( .A(n128), .B(n129), .Z(n131) );
  GTECH_XOR3 U112 ( .A(n132), .B(n122), .C(n121), .Z(n127) );
  GTECH_XOR2 U113 ( .A(n133), .B(n124), .Z(n121) );
  GTECH_OA22 U114 ( .A(n134), .B(n135), .C(n136), .D(n137), .Z(n124) );
  GTECH_NOR2 U115 ( .A(n138), .B(n139), .Z(n136) );
  GTECH_OR_NOT U116 ( .A(n140), .B(I_a[7]), .Z(n133) );
  GTECH_NOT U117 ( .A(n123), .Z(n122) );
  GTECH_XOR3 U118 ( .A(n115), .B(n114), .C(n116), .Z(n123) );
  GTECH_OAI21 U119 ( .A(n141), .B(n142), .C(n143), .Z(n116) );
  GTECH_OAI21 U120 ( .A(n144), .B(n145), .C(n146), .Z(n143) );
  GTECH_NOT U121 ( .A(n112), .Z(n114) );
  GTECH_OR_NOT U122 ( .A(n118), .B(I_b[6]), .Z(n112) );
  GTECH_NOT U123 ( .A(I_a[6]), .Z(n118) );
  GTECH_NOT U124 ( .A(n111), .Z(n115) );
  GTECH_OR_NOT U125 ( .A(n147), .B(I_b[7]), .Z(n111) );
  GTECH_NOT U126 ( .A(n119), .Z(n132) );
  GTECH_AO22 U127 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n119) );
  GTECH_OR2 U128 ( .A(n151), .B(n150), .Z(n149) );
  GTECH_XOR3 U129 ( .A(n152), .B(n153), .C(n128), .Z(N151) );
  GTECH_XOR3 U130 ( .A(n154), .B(n155), .C(n150), .Z(n128) );
  GTECH_XOR3 U131 ( .A(n134), .B(n135), .C(n137), .Z(n150) );
  GTECH_OAI21 U132 ( .A(n156), .B(n157), .C(n158), .Z(n137) );
  GTECH_OAI21 U133 ( .A(n159), .B(n160), .C(n161), .Z(n158) );
  GTECH_NOT U134 ( .A(n139), .Z(n135) );
  GTECH_OR_NOT U135 ( .A(n162), .B(I_a[7]), .Z(n139) );
  GTECH_NOT U136 ( .A(n138), .Z(n134) );
  GTECH_OR_NOT U137 ( .A(n140), .B(I_a[6]), .Z(n138) );
  GTECH_NOT U138 ( .A(I_b[5]), .Z(n140) );
  GTECH_NOT U139 ( .A(n151), .Z(n155) );
  GTECH_XOR3 U140 ( .A(n145), .B(n144), .C(n146), .Z(n151) );
  GTECH_OAI21 U141 ( .A(n163), .B(n164), .C(n165), .Z(n146) );
  GTECH_OAI21 U142 ( .A(n166), .B(n167), .C(n168), .Z(n165) );
  GTECH_NOT U143 ( .A(n142), .Z(n144) );
  GTECH_OR_NOT U144 ( .A(n147), .B(I_b[6]), .Z(n142) );
  GTECH_NOT U145 ( .A(n141), .Z(n145) );
  GTECH_OR_NOT U146 ( .A(n169), .B(I_b[7]), .Z(n141) );
  GTECH_NOT U147 ( .A(n148), .Z(n154) );
  GTECH_AO22 U148 ( .A(n170), .B(n171), .C(n172), .D(n173), .Z(n148) );
  GTECH_OR2 U149 ( .A(n173), .B(n172), .Z(n171) );
  GTECH_NOT U150 ( .A(n129), .Z(n153) );
  GTECH_OAI22 U151 ( .A(n174), .B(n175), .C(n105), .D(n176), .Z(n129) );
  GTECH_NOT U152 ( .A(n130), .Z(n152) );
  GTECH_AO22 U153 ( .A(n177), .B(n178), .C(n179), .D(n180), .Z(n130) );
  GTECH_OR2 U154 ( .A(n180), .B(n179), .Z(n178) );
  GTECH_XOR3 U155 ( .A(n181), .B(n182), .C(n179), .Z(N150) );
  GTECH_XOR3 U156 ( .A(n183), .B(n184), .C(n172), .Z(n179) );
  GTECH_XOR3 U157 ( .A(n160), .B(n159), .C(n161), .Z(n172) );
  GTECH_OAI21 U158 ( .A(n185), .B(n186), .C(n187), .Z(n161) );
  GTECH_OAI21 U159 ( .A(n188), .B(n189), .C(n190), .Z(n187) );
  GTECH_NOT U160 ( .A(n157), .Z(n159) );
  GTECH_OR_NOT U161 ( .A(n162), .B(I_a[6]), .Z(n157) );
  GTECH_NOT U162 ( .A(n156), .Z(n160) );
  GTECH_OR_NOT U163 ( .A(n147), .B(I_b[5]), .Z(n156) );
  GTECH_NOT U164 ( .A(I_a[5]), .Z(n147) );
  GTECH_NOT U165 ( .A(n173), .Z(n184) );
  GTECH_XOR3 U166 ( .A(n167), .B(n166), .C(n168), .Z(n173) );
  GTECH_OAI21 U167 ( .A(n191), .B(n192), .C(n193), .Z(n168) );
  GTECH_OAI21 U168 ( .A(n194), .B(n195), .C(n196), .Z(n193) );
  GTECH_NOT U169 ( .A(n164), .Z(n166) );
  GTECH_OR_NOT U170 ( .A(n169), .B(I_b[6]), .Z(n164) );
  GTECH_NOT U171 ( .A(n163), .Z(n167) );
  GTECH_OR_NOT U172 ( .A(n197), .B(I_b[7]), .Z(n163) );
  GTECH_NOT U173 ( .A(n170), .Z(n183) );
  GTECH_AO22 U174 ( .A(n198), .B(n199), .C(n200), .D(n201), .Z(n170) );
  GTECH_OR2 U175 ( .A(n201), .B(n200), .Z(n199) );
  GTECH_NOT U176 ( .A(n180), .Z(n182) );
  GTECH_XOR2 U177 ( .A(n175), .B(n174), .Z(n180) );
  GTECH_AND2 U178 ( .A(n202), .B(n203), .Z(n174) );
  GTECH_OR_NOT U179 ( .A(n204), .B(n205), .Z(n203) );
  GTECH_OAI21 U180 ( .A(n206), .B(n205), .C(n207), .Z(n202) );
  GTECH_XOR2 U181 ( .A(n208), .B(n176), .Z(n175) );
  GTECH_OAI22 U182 ( .A(n209), .B(n210), .C(n211), .D(n212), .Z(n176) );
  GTECH_NOR2 U183 ( .A(n213), .B(n214), .Z(n209) );
  GTECH_AND2 U184 ( .A(I_b[3]), .B(I_a[7]), .Z(n208) );
  GTECH_NOT U185 ( .A(n177), .Z(n181) );
  GTECH_OAI21 U186 ( .A(n215), .B(n216), .C(n217), .Z(n177) );
  GTECH_OAI21 U187 ( .A(n218), .B(n219), .C(n220), .Z(n217) );
  GTECH_XOR3 U188 ( .A(n221), .B(n216), .C(n219), .Z(N149) );
  GTECH_NOT U189 ( .A(n215), .Z(n219) );
  GTECH_XOR3 U190 ( .A(n206), .B(n222), .C(n205), .Z(n215) );
  GTECH_XOR3 U191 ( .A(n211), .B(n212), .C(n210), .Z(n205) );
  GTECH_OAI21 U192 ( .A(n223), .B(n224), .C(n225), .Z(n210) );
  GTECH_OAI21 U193 ( .A(n226), .B(n227), .C(n228), .Z(n225) );
  GTECH_NOT U194 ( .A(n214), .Z(n212) );
  GTECH_OR_NOT U195 ( .A(n229), .B(I_a[7]), .Z(n214) );
  GTECH_NOT U196 ( .A(n213), .Z(n211) );
  GTECH_OR_NOT U197 ( .A(n230), .B(I_a[6]), .Z(n213) );
  GTECH_NOT U198 ( .A(n207), .Z(n222) );
  GTECH_OAI2N2 U199 ( .A(n231), .B(n232), .C(n233), .D(n234), .Z(n207) );
  GTECH_OR_NOT U200 ( .A(n235), .B(n231), .Z(n234) );
  GTECH_NOT U201 ( .A(n204), .Z(n206) );
  GTECH_OR_NOT U202 ( .A(n105), .B(n236), .Z(n204) );
  GTECH_NOT U203 ( .A(I_a[7]), .Z(n105) );
  GTECH_NOT U204 ( .A(n218), .Z(n216) );
  GTECH_XOR3 U205 ( .A(n237), .B(n238), .C(n200), .Z(n218) );
  GTECH_XOR3 U206 ( .A(n189), .B(n188), .C(n190), .Z(n200) );
  GTECH_OAI21 U207 ( .A(n239), .B(n240), .C(n241), .Z(n190) );
  GTECH_OAI21 U208 ( .A(n242), .B(n243), .C(n244), .Z(n241) );
  GTECH_NOT U209 ( .A(n186), .Z(n188) );
  GTECH_OR_NOT U210 ( .A(n162), .B(I_a[5]), .Z(n186) );
  GTECH_NOT U211 ( .A(I_b[4]), .Z(n162) );
  GTECH_NOT U212 ( .A(n185), .Z(n189) );
  GTECH_OR_NOT U213 ( .A(n169), .B(I_b[5]), .Z(n185) );
  GTECH_NOT U214 ( .A(n201), .Z(n238) );
  GTECH_XOR3 U215 ( .A(n195), .B(n194), .C(n196), .Z(n201) );
  GTECH_OAI21 U216 ( .A(n245), .B(n246), .C(n247), .Z(n196) );
  GTECH_NOT U217 ( .A(n192), .Z(n194) );
  GTECH_OR_NOT U218 ( .A(n197), .B(I_b[6]), .Z(n192) );
  GTECH_NOT U219 ( .A(n191), .Z(n195) );
  GTECH_OR_NOT U220 ( .A(n248), .B(I_b[7]), .Z(n191) );
  GTECH_NOT U221 ( .A(n198), .Z(n237) );
  GTECH_OAI2N2 U222 ( .A(n249), .B(n250), .C(n251), .D(n252), .Z(n198) );
  GTECH_OR_NOT U223 ( .A(n253), .B(n249), .Z(n252) );
  GTECH_NOT U224 ( .A(n220), .Z(n221) );
  GTECH_OAI2N2 U225 ( .A(n254), .B(n255), .C(n256), .D(n257), .Z(n220) );
  GTECH_OR_NOT U226 ( .A(n258), .B(n254), .Z(n257) );
  GTECH_XOR3 U227 ( .A(n259), .B(n258), .C(n254), .Z(N148) );
  GTECH_XOR3 U228 ( .A(n260), .B(n232), .C(n231), .Z(n254) );
  GTECH_XOR2 U229 ( .A(n261), .B(n236), .Z(n231) );
  GTECH_OA21 U230 ( .A(n262), .B(n263), .C(n264), .Z(n236) );
  GTECH_OAI21 U231 ( .A(n265), .B(n266), .C(n267), .Z(n264) );
  GTECH_OR_NOT U232 ( .A(n268), .B(I_a[7]), .Z(n261) );
  GTECH_NOT U233 ( .A(n235), .Z(n232) );
  GTECH_XOR3 U234 ( .A(n227), .B(n226), .C(n228), .Z(n235) );
  GTECH_OAI21 U235 ( .A(n269), .B(n270), .C(n271), .Z(n228) );
  GTECH_OAI21 U236 ( .A(n272), .B(n273), .C(n274), .Z(n271) );
  GTECH_NOT U237 ( .A(n224), .Z(n226) );
  GTECH_OR_NOT U238 ( .A(n229), .B(I_a[6]), .Z(n224) );
  GTECH_NOT U239 ( .A(n223), .Z(n227) );
  GTECH_OR_NOT U240 ( .A(n230), .B(I_a[5]), .Z(n223) );
  GTECH_NOT U241 ( .A(n233), .Z(n260) );
  GTECH_OAI2N2 U242 ( .A(n275), .B(n276), .C(n277), .D(n278), .Z(n233) );
  GTECH_OR_NOT U243 ( .A(n279), .B(n275), .Z(n278) );
  GTECH_NOT U244 ( .A(n255), .Z(n258) );
  GTECH_XOR3 U245 ( .A(n280), .B(n250), .C(n249), .Z(n255) );
  GTECH_XOR3 U246 ( .A(n281), .B(n282), .C(n247), .Z(n249) );
  GTECH_NAND3 U247 ( .A(I_b[6]), .B(I_a[1]), .C(n283), .Z(n247) );
  GTECH_NOT U248 ( .A(n246), .Z(n282) );
  GTECH_OR_NOT U249 ( .A(n248), .B(I_b[6]), .Z(n246) );
  GTECH_NOT U250 ( .A(n245), .Z(n281) );
  GTECH_OR_NOT U251 ( .A(n284), .B(I_b[7]), .Z(n245) );
  GTECH_NOT U252 ( .A(n253), .Z(n250) );
  GTECH_XOR3 U253 ( .A(n243), .B(n242), .C(n244), .Z(n253) );
  GTECH_OAI21 U254 ( .A(n285), .B(n286), .C(n287), .Z(n244) );
  GTECH_OAI21 U255 ( .A(n288), .B(n289), .C(n290), .Z(n287) );
  GTECH_NOT U256 ( .A(n240), .Z(n242) );
  GTECH_OR_NOT U257 ( .A(n169), .B(I_b[4]), .Z(n240) );
  GTECH_NOT U258 ( .A(I_a[4]), .Z(n169) );
  GTECH_NOT U259 ( .A(n239), .Z(n243) );
  GTECH_OR_NOT U260 ( .A(n197), .B(I_b[5]), .Z(n239) );
  GTECH_NOT U261 ( .A(n251), .Z(n280) );
  GTECH_OAI22 U262 ( .A(n291), .B(n292), .C(n293), .D(n294), .Z(n251) );
  GTECH_AND_NOT U263 ( .A(n293), .B(n295), .Z(n291) );
  GTECH_NOT U264 ( .A(n256), .Z(n259) );
  GTECH_OAI21 U265 ( .A(n296), .B(n297), .C(n298), .Z(n256) );
  GTECH_OAI21 U266 ( .A(n299), .B(n300), .C(n301), .Z(n298) );
  GTECH_XOR3 U267 ( .A(n302), .B(n297), .C(n300), .Z(N147) );
  GTECH_NOT U268 ( .A(n296), .Z(n300) );
  GTECH_XOR3 U269 ( .A(n303), .B(n276), .C(n275), .Z(n296) );
  GTECH_XOR3 U270 ( .A(n262), .B(n263), .C(n267), .Z(n275) );
  GTECH_OAI21 U271 ( .A(n304), .B(n305), .C(n306), .Z(n267) );
  GTECH_OAI21 U272 ( .A(n307), .B(n308), .C(n309), .Z(n306) );
  GTECH_NOT U273 ( .A(n266), .Z(n263) );
  GTECH_OR_NOT U274 ( .A(n310), .B(I_a[7]), .Z(n266) );
  GTECH_NOT U275 ( .A(n265), .Z(n262) );
  GTECH_OR_NOT U276 ( .A(n268), .B(I_a[6]), .Z(n265) );
  GTECH_NOT U277 ( .A(n279), .Z(n276) );
  GTECH_XOR3 U278 ( .A(n273), .B(n272), .C(n274), .Z(n279) );
  GTECH_OAI21 U279 ( .A(n311), .B(n312), .C(n313), .Z(n274) );
  GTECH_OAI21 U280 ( .A(n314), .B(n315), .C(n316), .Z(n313) );
  GTECH_NOT U281 ( .A(n270), .Z(n272) );
  GTECH_OR_NOT U282 ( .A(n229), .B(I_a[5]), .Z(n270) );
  GTECH_NOT U283 ( .A(n269), .Z(n273) );
  GTECH_OR_NOT U284 ( .A(n230), .B(I_a[4]), .Z(n269) );
  GTECH_NOT U285 ( .A(n277), .Z(n303) );
  GTECH_OAI2N2 U286 ( .A(n317), .B(n318), .C(n319), .D(n320), .Z(n277) );
  GTECH_OR_NOT U287 ( .A(n321), .B(n317), .Z(n320) );
  GTECH_NOT U288 ( .A(n299), .Z(n297) );
  GTECH_XOR3 U289 ( .A(n322), .B(n294), .C(n293), .Z(n299) );
  GTECH_XOR2 U290 ( .A(n323), .B(n283), .Z(n293) );
  GTECH_NOT U291 ( .A(n324), .Z(n283) );
  GTECH_OR_NOT U292 ( .A(n325), .B(I_b[7]), .Z(n324) );
  GTECH_OR_NOT U293 ( .A(n284), .B(I_b[6]), .Z(n323) );
  GTECH_NOT U294 ( .A(n295), .Z(n294) );
  GTECH_XOR3 U295 ( .A(n289), .B(n288), .C(n290), .Z(n295) );
  GTECH_OAI21 U296 ( .A(n326), .B(n327), .C(n328), .Z(n290) );
  GTECH_NOT U297 ( .A(n286), .Z(n288) );
  GTECH_OR_NOT U298 ( .A(n197), .B(I_b[4]), .Z(n286) );
  GTECH_NOT U299 ( .A(I_a[3]), .Z(n197) );
  GTECH_NOT U300 ( .A(n285), .Z(n289) );
  GTECH_OR_NOT U301 ( .A(n248), .B(I_b[5]), .Z(n285) );
  GTECH_NOT U302 ( .A(n292), .Z(n322) );
  GTECH_NAND3 U303 ( .A(I_a[0]), .B(n329), .C(I_b[6]), .Z(n292) );
  GTECH_NOT U304 ( .A(n330), .Z(n329) );
  GTECH_NOT U305 ( .A(n301), .Z(n302) );
  GTECH_OAI2N2 U306 ( .A(n331), .B(n332), .C(n333), .D(n334), .Z(n301) );
  GTECH_OR_NOT U307 ( .A(n335), .B(n331), .Z(n334) );
  GTECH_XOR3 U308 ( .A(n336), .B(n335), .C(n331), .Z(N146) );
  GTECH_XOR3 U309 ( .A(n337), .B(n318), .C(n317), .Z(n331) );
  GTECH_XOR3 U310 ( .A(n304), .B(n305), .C(n309), .Z(n317) );
  GTECH_OAI21 U311 ( .A(n338), .B(n339), .C(n340), .Z(n309) );
  GTECH_OAI21 U312 ( .A(n341), .B(n342), .C(n343), .Z(n340) );
  GTECH_NOT U313 ( .A(n308), .Z(n305) );
  GTECH_OR_NOT U314 ( .A(n310), .B(I_a[6]), .Z(n308) );
  GTECH_NOT U315 ( .A(n307), .Z(n304) );
  GTECH_OR_NOT U316 ( .A(n268), .B(I_a[5]), .Z(n307) );
  GTECH_NOT U317 ( .A(n321), .Z(n318) );
  GTECH_XOR3 U318 ( .A(n315), .B(n314), .C(n316), .Z(n321) );
  GTECH_OAI21 U319 ( .A(n344), .B(n345), .C(n346), .Z(n316) );
  GTECH_OAI21 U320 ( .A(n347), .B(n348), .C(n349), .Z(n346) );
  GTECH_NOT U321 ( .A(n312), .Z(n314) );
  GTECH_OR_NOT U322 ( .A(n229), .B(I_a[4]), .Z(n312) );
  GTECH_NOT U323 ( .A(n311), .Z(n315) );
  GTECH_OR_NOT U324 ( .A(n230), .B(I_a[3]), .Z(n311) );
  GTECH_NOT U325 ( .A(n319), .Z(n337) );
  GTECH_OAI2N2 U326 ( .A(n350), .B(n351), .C(n352), .D(n353), .Z(n319) );
  GTECH_OR_NOT U327 ( .A(n354), .B(n350), .Z(n353) );
  GTECH_NOT U328 ( .A(n332), .Z(n335) );
  GTECH_XOR2 U329 ( .A(n330), .B(n355), .Z(n332) );
  GTECH_AND2 U330 ( .A(I_b[6]), .B(I_a[0]), .Z(n355) );
  GTECH_XOR3 U331 ( .A(n356), .B(n357), .C(n328), .Z(n330) );
  GTECH_NAND3 U332 ( .A(I_b[4]), .B(I_a[1]), .C(n358), .Z(n328) );
  GTECH_NOT U333 ( .A(n327), .Z(n357) );
  GTECH_OR_NOT U334 ( .A(n248), .B(I_b[4]), .Z(n327) );
  GTECH_NOT U335 ( .A(n326), .Z(n356) );
  GTECH_OR_NOT U336 ( .A(n284), .B(I_b[5]), .Z(n326) );
  GTECH_NOT U337 ( .A(n333), .Z(n336) );
  GTECH_OAI21 U338 ( .A(n359), .B(n360), .C(n361), .Z(n333) );
  GTECH_OAI21 U339 ( .A(n362), .B(n363), .C(n364), .Z(n361) );
  GTECH_XOR3 U340 ( .A(n364), .B(n362), .C(n363), .Z(N145) );
  GTECH_NOT U341 ( .A(n359), .Z(n363) );
  GTECH_XOR3 U342 ( .A(n365), .B(n351), .C(n350), .Z(n359) );
  GTECH_XOR3 U343 ( .A(n338), .B(n339), .C(n343), .Z(n350) );
  GTECH_OAI21 U344 ( .A(n366), .B(n367), .C(n368), .Z(n343) );
  GTECH_OAI21 U345 ( .A(n369), .B(n370), .C(n371), .Z(n368) );
  GTECH_NOT U346 ( .A(n342), .Z(n339) );
  GTECH_OR_NOT U347 ( .A(n310), .B(I_a[5]), .Z(n342) );
  GTECH_NOT U348 ( .A(n341), .Z(n338) );
  GTECH_OR_NOT U349 ( .A(n268), .B(I_a[4]), .Z(n341) );
  GTECH_NOT U350 ( .A(n354), .Z(n351) );
  GTECH_XOR3 U351 ( .A(n348), .B(n347), .C(n349), .Z(n354) );
  GTECH_OAI21 U352 ( .A(n372), .B(n373), .C(n374), .Z(n349) );
  GTECH_NOT U353 ( .A(n345), .Z(n347) );
  GTECH_OR_NOT U354 ( .A(n229), .B(I_a[3]), .Z(n345) );
  GTECH_NOT U355 ( .A(n344), .Z(n348) );
  GTECH_OR_NOT U356 ( .A(n230), .B(I_a[2]), .Z(n344) );
  GTECH_NOT U357 ( .A(n352), .Z(n365) );
  GTECH_OAI2N2 U358 ( .A(n375), .B(n376), .C(n377), .D(n378), .Z(n352) );
  GTECH_OR_NOT U359 ( .A(n379), .B(n375), .Z(n378) );
  GTECH_NOT U360 ( .A(n360), .Z(n362) );
  GTECH_XOR2 U361 ( .A(n380), .B(n358), .Z(n360) );
  GTECH_NOT U362 ( .A(n381), .Z(n358) );
  GTECH_OR_NOT U363 ( .A(n325), .B(I_b[5]), .Z(n381) );
  GTECH_OR_NOT U364 ( .A(n284), .B(I_b[4]), .Z(n380) );
  GTECH_NOT U365 ( .A(n382), .Z(n364) );
  GTECH_NAND3 U366 ( .A(n383), .B(I_a[0]), .C(I_b[4]), .Z(n382) );
  GTECH_XOR2 U367 ( .A(n383), .B(n384), .Z(N144) );
  GTECH_AND2 U368 ( .A(I_b[4]), .B(I_a[0]), .Z(n384) );
  GTECH_XOR3 U369 ( .A(n385), .B(n379), .C(n375), .Z(n383) );
  GTECH_XOR3 U370 ( .A(n386), .B(n387), .C(n374), .Z(n375) );
  GTECH_NAND3 U371 ( .A(I_a[1]), .B(n388), .C(I_b[2]), .Z(n374) );
  GTECH_NOT U372 ( .A(n373), .Z(n387) );
  GTECH_OR_NOT U373 ( .A(n229), .B(I_a[2]), .Z(n373) );
  GTECH_NOT U374 ( .A(I_b[2]), .Z(n229) );
  GTECH_NOT U375 ( .A(n372), .Z(n386) );
  GTECH_OR_NOT U376 ( .A(n230), .B(I_a[1]), .Z(n372) );
  GTECH_NOT U377 ( .A(I_b[3]), .Z(n230) );
  GTECH_NOT U378 ( .A(n376), .Z(n379) );
  GTECH_XOR3 U379 ( .A(n366), .B(n367), .C(n371), .Z(n376) );
  GTECH_OAI22 U380 ( .A(n389), .B(n390), .C(n391), .D(n392), .Z(n371) );
  GTECH_NOR2 U381 ( .A(n393), .B(n394), .Z(n389) );
  GTECH_NOT U382 ( .A(n370), .Z(n367) );
  GTECH_OR_NOT U383 ( .A(n310), .B(I_a[4]), .Z(n370) );
  GTECH_NOT U384 ( .A(n369), .Z(n366) );
  GTECH_OR_NOT U385 ( .A(n268), .B(I_a[3]), .Z(n369) );
  GTECH_NOT U386 ( .A(I_b[1]), .Z(n268) );
  GTECH_NOT U387 ( .A(n377), .Z(n385) );
  GTECH_OAI21 U388 ( .A(n395), .B(n396), .C(n397), .Z(n377) );
  GTECH_OAI21 U389 ( .A(n398), .B(n399), .C(n400), .Z(n397) );
  GTECH_NOT U390 ( .A(n399), .Z(n395) );
  GTECH_XOR3 U391 ( .A(n400), .B(n398), .C(n399), .Z(N143) );
  GTECH_XOR3 U392 ( .A(n391), .B(n392), .C(n390), .Z(n399) );
  GTECH_OAI21 U393 ( .A(n401), .B(n402), .C(n403), .Z(n390) );
  GTECH_NOT U394 ( .A(n394), .Z(n392) );
  GTECH_OR_NOT U395 ( .A(n310), .B(I_a[3]), .Z(n394) );
  GTECH_NOT U396 ( .A(I_b[0]), .Z(n310) );
  GTECH_NOT U397 ( .A(n393), .Z(n391) );
  GTECH_OR_NOT U398 ( .A(n248), .B(I_b[1]), .Z(n393) );
  GTECH_NOT U399 ( .A(n396), .Z(n398) );
  GTECH_XOR2 U400 ( .A(n404), .B(n388), .Z(n396) );
  GTECH_NOT U401 ( .A(n405), .Z(n388) );
  GTECH_OR_NOT U402 ( .A(n325), .B(I_b[3]), .Z(n405) );
  GTECH_OR_NOT U403 ( .A(n284), .B(I_b[2]), .Z(n404) );
  GTECH_NOT U404 ( .A(n406), .Z(n400) );
  GTECH_NAND3 U405 ( .A(I_a[0]), .B(n407), .C(I_b[2]), .Z(n406) );
  GTECH_XOR2 U406 ( .A(n408), .B(n407), .Z(N142) );
  GTECH_NOT U407 ( .A(n409), .Z(n407) );
  GTECH_XOR3 U408 ( .A(n410), .B(n411), .C(n403), .Z(n409) );
  GTECH_NAND3 U409 ( .A(n412), .B(I_a[1]), .C(I_b[0]), .Z(n403) );
  GTECH_NOT U410 ( .A(n402), .Z(n411) );
  GTECH_OR_NOT U411 ( .A(n248), .B(I_b[0]), .Z(n402) );
  GTECH_NOT U412 ( .A(I_a[2]), .Z(n248) );
  GTECH_NOT U413 ( .A(n401), .Z(n410) );
  GTECH_OR_NOT U414 ( .A(n284), .B(I_b[1]), .Z(n401) );
  GTECH_NOT U415 ( .A(I_a[1]), .Z(n284) );
  GTECH_AND2 U416 ( .A(I_b[2]), .B(I_a[0]), .Z(n408) );
  GTECH_XOR2 U417 ( .A(n412), .B(n413), .Z(N141) );
  GTECH_AND2 U418 ( .A(I_b[0]), .B(I_a[1]), .Z(n413) );
  GTECH_NOT U419 ( .A(n414), .Z(n412) );
  GTECH_OR_NOT U420 ( .A(n325), .B(I_b[1]), .Z(n414) );
  GTECH_NOT U421 ( .A(I_a[0]), .Z(n325) );
  GTECH_AND2 U422 ( .A(I_b[0]), .B(I_a[0]), .Z(N140) );
endmodule

