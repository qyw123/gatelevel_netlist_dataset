
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169;

  GTECH_XNOR2 U103 ( .A(n84), .B(n85), .Z(sum[9]) );
  GTECH_XOR2 U104 ( .A(n86), .B(n87), .Z(sum[8]) );
  GTECH_XOR2 U105 ( .A(n88), .B(n89), .Z(sum[7]) );
  GTECH_AO21 U106 ( .A(n90), .B(n91), .C(n92), .Z(n88) );
  GTECH_XOR2 U107 ( .A(n90), .B(n91), .Z(sum[6]) );
  GTECH_AO21 U108 ( .A(n93), .B(n94), .C(n95), .Z(n90) );
  GTECH_XOR2 U109 ( .A(n94), .B(n93), .Z(sum[5]) );
  GTECH_AO21 U110 ( .A(n96), .B(n97), .C(n98), .Z(n93) );
  GTECH_XOR2 U111 ( .A(n97), .B(n96), .Z(sum[4]) );
  GTECH_XNOR2 U112 ( .A(n99), .B(n100), .Z(sum[3]) );
  GTECH_AOI21 U113 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_XOR2 U114 ( .A(n101), .B(n102), .Z(sum[2]) );
  GTECH_AO21 U115 ( .A(n104), .B(n105), .C(n106), .Z(n101) );
  GTECH_XOR2 U116 ( .A(n104), .B(n105), .Z(sum[1]) );
  GTECH_NOT U117 ( .A(n107), .Z(n104) );
  GTECH_AOI22 U118 ( .A(a[0]), .B(b[0]), .C(n108), .D(cin), .Z(n107) );
  GTECH_XOR2 U119 ( .A(n109), .B(n110), .Z(sum[15]) );
  GTECH_OA21 U120 ( .A(n111), .B(n112), .C(n113), .Z(n110) );
  GTECH_XOR2 U121 ( .A(n111), .B(n112), .Z(sum[14]) );
  GTECH_AOI21 U122 ( .A(n114), .B(n115), .C(n116), .Z(n111) );
  GTECH_NOT U123 ( .A(n117), .Z(n115) );
  GTECH_XNOR2 U124 ( .A(n117), .B(n114), .Z(sum[13]) );
  GTECH_AO21 U125 ( .A(cout), .B(n118), .C(n119), .Z(n114) );
  GTECH_XNOR2 U126 ( .A(cout), .B(n120), .Z(sum[12]) );
  GTECH_XNOR2 U127 ( .A(n121), .B(n122), .Z(sum[11]) );
  GTECH_AO21 U128 ( .A(n123), .B(n124), .C(n125), .Z(n121) );
  GTECH_XNOR2 U129 ( .A(n126), .B(n123), .Z(sum[10]) );
  GTECH_OAI21 U130 ( .A(n84), .B(n127), .C(n128), .Z(n123) );
  GTECH_AOI2N2 U131 ( .A(a[8]), .B(b[8]), .C(n87), .D(n86), .Z(n84) );
  GTECH_XOR2 U132 ( .A(cin), .B(n108), .Z(sum[0]) );
  GTECH_OAI21 U133 ( .A(n87), .B(n129), .C(n130), .Z(cout) );
  GTECH_AOI21 U134 ( .A(n96), .B(n131), .C(n132), .Z(n87) );
  GTECH_OAI21 U135 ( .A(n133), .B(n134), .C(n135), .Z(n96) );
  GTECH_NAND3 U136 ( .A(n136), .B(n102), .C(cin), .Z(n134) );
  GTECH_NAND3 U137 ( .A(n108), .B(n99), .C(n105), .Z(n133) );
  GTECH_AND4 U138 ( .A(n131), .B(n136), .C(n137), .D(n138), .Z(Pm) );
  GTECH_AND4 U139 ( .A(n102), .B(n105), .C(n108), .D(n99), .Z(n138) );
  GTECH_XOR2 U140 ( .A(a[0]), .B(b[0]), .Z(n108) );
  GTECH_OAI21 U141 ( .A(n139), .B(n129), .C(n130), .Z(Gm) );
  GTECH_AOI2N2 U142 ( .A(b[15]), .B(a[15]), .C(n140), .D(n109), .Z(n130) );
  GTECH_OA21 U143 ( .A(n141), .B(n112), .C(n113), .Z(n140) );
  GTECH_OA21 U144 ( .A(n117), .B(n142), .C(n143), .Z(n141) );
  GTECH_NOT U145 ( .A(n137), .Z(n129) );
  GTECH_NOR4 U146 ( .A(n120), .B(n112), .C(n117), .D(n109), .Z(n137) );
  GTECH_XNOR2 U147 ( .A(a[15]), .B(b[15]), .Z(n109) );
  GTECH_OAI21 U148 ( .A(b[13]), .B(a[13]), .C(n143), .Z(n117) );
  GTECH_NOT U149 ( .A(n116), .Z(n143) );
  GTECH_AND2 U150 ( .A(b[13]), .B(a[13]), .Z(n116) );
  GTECH_OAI21 U151 ( .A(a[14]), .B(b[14]), .C(n113), .Z(n112) );
  GTECH_NOT U152 ( .A(n144), .Z(n113) );
  GTECH_AND2 U153 ( .A(a[14]), .B(b[14]), .Z(n144) );
  GTECH_NOT U154 ( .A(n118), .Z(n120) );
  GTECH_OA21 U155 ( .A(b[12]), .B(a[12]), .C(n142), .Z(n118) );
  GTECH_NOT U156 ( .A(n119), .Z(n142) );
  GTECH_AND2 U157 ( .A(b[12]), .B(a[12]), .Z(n119) );
  GTECH_AOI21 U158 ( .A(n145), .B(n131), .C(n132), .Z(n139) );
  GTECH_OAI21 U159 ( .A(n146), .B(n122), .C(n147), .Z(n132) );
  GTECH_AND2 U160 ( .A(n148), .B(n149), .Z(n146) );
  GTECH_OAI21 U161 ( .A(n150), .B(n151), .C(n124), .Z(n148) );
  GTECH_AND3 U162 ( .A(a[8]), .B(n85), .C(b[8]), .Z(n151) );
  GTECH_NOR4 U163 ( .A(n122), .B(n126), .C(n127), .D(n86), .Z(n131) );
  GTECH_XNOR2 U164 ( .A(a[8]), .B(b[8]), .Z(n86) );
  GTECH_NOT U165 ( .A(n85), .Z(n127) );
  GTECH_OA21 U166 ( .A(a[9]), .B(b[9]), .C(n128), .Z(n85) );
  GTECH_NOT U167 ( .A(n150), .Z(n128) );
  GTECH_AND2 U168 ( .A(b[9]), .B(a[9]), .Z(n150) );
  GTECH_NOT U169 ( .A(n124), .Z(n126) );
  GTECH_OA21 U170 ( .A(b[10]), .B(a[10]), .C(n149), .Z(n124) );
  GTECH_NOT U171 ( .A(n125), .Z(n149) );
  GTECH_AND2 U172 ( .A(a[10]), .B(b[10]), .Z(n125) );
  GTECH_OAI21 U173 ( .A(b[11]), .B(a[11]), .C(n147), .Z(n122) );
  GTECH_OR_NOT U174 ( .A(n152), .B(a[11]), .Z(n147) );
  GTECH_NOT U175 ( .A(b[11]), .Z(n152) );
  GTECH_NOT U176 ( .A(n135), .Z(n145) );
  GTECH_OA21 U177 ( .A(n153), .B(n154), .C(n155), .Z(n135) );
  GTECH_AOI21 U178 ( .A(n156), .B(n136), .C(n157), .Z(n155) );
  GTECH_AND4 U179 ( .A(n91), .B(n97), .C(n89), .D(n94), .Z(n136) );
  GTECH_OA21 U180 ( .A(b[4]), .B(a[4]), .C(n158), .Z(n97) );
  GTECH_NOT U181 ( .A(n98), .Z(n158) );
  GTECH_AO21 U182 ( .A(b[3]), .B(a[3]), .C(n159), .Z(n156) );
  GTECH_NOT U183 ( .A(n160), .Z(n159) );
  GTECH_OAI21 U184 ( .A(n103), .B(n161), .C(n99), .Z(n160) );
  GTECH_XNOR2 U185 ( .A(a[3]), .B(n162), .Z(n99) );
  GTECH_NOT U186 ( .A(b[3]), .Z(n162) );
  GTECH_OA21 U187 ( .A(n106), .B(n163), .C(n102), .Z(n161) );
  GTECH_OA21 U188 ( .A(a[2]), .B(b[2]), .C(n164), .Z(n102) );
  GTECH_NOT U189 ( .A(n103), .Z(n164) );
  GTECH_AND3 U190 ( .A(a[0]), .B(n105), .C(b[0]), .Z(n163) );
  GTECH_OA21 U191 ( .A(a[1]), .B(b[1]), .C(n165), .Z(n105) );
  GTECH_NOT U192 ( .A(n106), .Z(n165) );
  GTECH_AND2 U193 ( .A(b[1]), .B(a[1]), .Z(n106) );
  GTECH_AND2 U194 ( .A(b[2]), .B(a[2]), .Z(n103) );
  GTECH_NOT U195 ( .A(n89), .Z(n154) );
  GTECH_OA21 U196 ( .A(b[7]), .B(a[7]), .C(n166), .Z(n89) );
  GTECH_NOT U197 ( .A(n157), .Z(n166) );
  GTECH_AND2 U198 ( .A(b[7]), .B(a[7]), .Z(n157) );
  GTECH_AOI21 U199 ( .A(n167), .B(n91), .C(n92), .Z(n153) );
  GTECH_OA21 U200 ( .A(a[6]), .B(b[6]), .C(n168), .Z(n91) );
  GTECH_NOT U201 ( .A(n92), .Z(n168) );
  GTECH_AND2 U202 ( .A(a[6]), .B(b[6]), .Z(n92) );
  GTECH_AO21 U203 ( .A(n94), .B(n98), .C(n95), .Z(n167) );
  GTECH_AND2 U204 ( .A(b[4]), .B(a[4]), .Z(n98) );
  GTECH_OA21 U205 ( .A(b[5]), .B(a[5]), .C(n169), .Z(n94) );
  GTECH_NOT U206 ( .A(n95), .Z(n169) );
  GTECH_AND2 U207 ( .A(b[5]), .B(a[5]), .Z(n95) );
endmodule

