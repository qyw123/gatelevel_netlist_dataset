
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NAND2 U83 ( .A(n93), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI22 U86 ( .A(n98), .B(n99), .C(n100), .D(n101), .Z(n89) );
  GTECH_AND_NOT U87 ( .A(n98), .B(n102), .Z(n100) );
  GTECH_NOT U88 ( .A(n103), .Z(n98) );
  GTECH_NAND2 U89 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n104), .Z(n84) );
  GTECH_NAND2 U91 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_XOR2 U92 ( .A(n106), .B(n105), .Z(N153) );
  GTECH_NOT U93 ( .A(n107), .Z(n105) );
  GTECH_XOR3 U94 ( .A(n108), .B(n93), .C(n95), .Z(n107) );
  GTECH_XOR3 U95 ( .A(n102), .B(n109), .C(n103), .Z(n95) );
  GTECH_OAI22 U96 ( .A(n110), .B(n111), .C(n112), .D(n113), .Z(n103) );
  GTECH_AND_NOT U97 ( .A(n110), .B(n114), .Z(n112) );
  GTECH_NOT U98 ( .A(n115), .Z(n110) );
  GTECH_NOT U99 ( .A(n101), .Z(n109) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n101) );
  GTECH_NOT U101 ( .A(n99), .Z(n102) );
  GTECH_NAND2 U102 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U103 ( .A(n116), .B(n117), .C(n118), .COUT(n93) );
  GTECH_NOT U104 ( .A(n119), .Z(n118) );
  GTECH_XOR2 U105 ( .A(n120), .B(n121), .Z(n117) );
  GTECH_AND_NOT U106 ( .A(I_a[7]), .B(n122), .Z(n121) );
  GTECH_NOT U107 ( .A(I_b[5]), .Z(n122) );
  GTECH_NOT U108 ( .A(n123), .Z(n120) );
  GTECH_NOT U109 ( .A(n94), .Z(n108) );
  GTECH_NAND2 U110 ( .A(I_a[7]), .B(n123), .Z(n94) );
  GTECH_NOT U111 ( .A(n124), .Z(n106) );
  GTECH_NAND2 U112 ( .A(n125), .B(n126), .Z(n124) );
  GTECH_NOT U113 ( .A(n127), .Z(n126) );
  GTECH_XOR2 U114 ( .A(n127), .B(n128), .Z(N152) );
  GTECH_NOT U115 ( .A(n125), .Z(n128) );
  GTECH_XOR4 U116 ( .A(n119), .B(n116), .C(n129), .D(n123), .Z(n125) );
  GTECH_OAI22 U117 ( .A(n130), .B(n131), .C(n132), .D(n133), .Z(n123) );
  GTECH_AND_NOT U118 ( .A(n130), .B(n134), .Z(n132) );
  GTECH_NAND2 U119 ( .A(I_a[7]), .B(I_b[5]), .Z(n129) );
  GTECH_ADD_ABC U120 ( .A(n135), .B(n136), .C(n137), .COUT(n116) );
  GTECH_NOT U121 ( .A(n138), .Z(n137) );
  GTECH_XOR3 U122 ( .A(n134), .B(n139), .C(n130), .Z(n136) );
  GTECH_NOT U123 ( .A(n140), .Z(n130) );
  GTECH_NOT U124 ( .A(n131), .Z(n134) );
  GTECH_XOR3 U125 ( .A(n114), .B(n141), .C(n115), .Z(n119) );
  GTECH_OAI22 U126 ( .A(n142), .B(n143), .C(n144), .D(n145), .Z(n115) );
  GTECH_AND_NOT U127 ( .A(n142), .B(n146), .Z(n144) );
  GTECH_NOT U128 ( .A(n147), .Z(n142) );
  GTECH_NOT U129 ( .A(n113), .Z(n141) );
  GTECH_NAND2 U130 ( .A(I_b[7]), .B(I_a[5]), .Z(n113) );
  GTECH_NOT U131 ( .A(n111), .Z(n114) );
  GTECH_NAND2 U132 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_ADD_ABC U133 ( .A(n148), .B(n149), .C(n150), .COUT(n127) );
  GTECH_NOT U134 ( .A(n151), .Z(n150) );
  GTECH_OA22 U135 ( .A(n152), .B(n153), .C(n154), .D(n155), .Z(n149) );
  GTECH_OA21 U136 ( .A(n156), .B(n157), .C(n158), .Z(n148) );
  GTECH_AO21 U137 ( .A(n156), .B(n157), .C(n159), .Z(n158) );
  GTECH_XOR3 U138 ( .A(n160), .B(n151), .C(n161), .Z(N151) );
  GTECH_OA21 U139 ( .A(n156), .B(n157), .C(n162), .Z(n161) );
  GTECH_AO21 U140 ( .A(n156), .B(n157), .C(n159), .Z(n162) );
  GTECH_XOR2 U141 ( .A(n163), .B(n135), .Z(n151) );
  GTECH_ADD_ABC U142 ( .A(n164), .B(n165), .C(n166), .COUT(n135) );
  GTECH_NOT U143 ( .A(n167), .Z(n166) );
  GTECH_XOR3 U144 ( .A(n168), .B(n169), .C(n170), .Z(n165) );
  GTECH_XOR4 U145 ( .A(n139), .B(n140), .C(n131), .D(n138), .Z(n163) );
  GTECH_XOR3 U146 ( .A(n146), .B(n171), .C(n147), .Z(n138) );
  GTECH_OAI22 U147 ( .A(n172), .B(n173), .C(n174), .D(n175), .Z(n147) );
  GTECH_AND_NOT U148 ( .A(n172), .B(n176), .Z(n174) );
  GTECH_NOT U149 ( .A(n177), .Z(n172) );
  GTECH_NOT U150 ( .A(n145), .Z(n171) );
  GTECH_NAND2 U151 ( .A(I_b[7]), .B(I_a[4]), .Z(n145) );
  GTECH_NOT U152 ( .A(n143), .Z(n146) );
  GTECH_NAND2 U153 ( .A(I_b[6]), .B(I_a[5]), .Z(n143) );
  GTECH_NAND2 U154 ( .A(I_a[7]), .B(I_b[4]), .Z(n131) );
  GTECH_OAI22 U155 ( .A(n170), .B(n178), .C(n179), .D(n180), .Z(n140) );
  GTECH_AND_NOT U156 ( .A(n170), .B(n168), .Z(n179) );
  GTECH_NOT U157 ( .A(n181), .Z(n170) );
  GTECH_NOT U158 ( .A(n133), .Z(n139) );
  GTECH_NAND2 U159 ( .A(I_a[6]), .B(I_b[5]), .Z(n133) );
  GTECH_OA22 U160 ( .A(n152), .B(n153), .C(n154), .D(n155), .Z(n160) );
  GTECH_NOT U161 ( .A(n182), .Z(n155) );
  GTECH_NOT U162 ( .A(I_a[7]), .Z(n153) );
  GTECH_XOR3 U163 ( .A(n156), .B(n183), .C(n159), .Z(N150) );
  GTECH_XOR2 U164 ( .A(n164), .B(n184), .Z(n159) );
  GTECH_XOR4 U165 ( .A(n169), .B(n181), .C(n167), .D(n168), .Z(n184) );
  GTECH_NOT U166 ( .A(n178), .Z(n168) );
  GTECH_NAND2 U167 ( .A(I_a[6]), .B(I_b[4]), .Z(n178) );
  GTECH_XOR3 U168 ( .A(n176), .B(n185), .C(n177), .Z(n167) );
  GTECH_OAI22 U169 ( .A(n186), .B(n187), .C(n188), .D(n189), .Z(n177) );
  GTECH_AND_NOT U170 ( .A(n186), .B(n190), .Z(n188) );
  GTECH_NOT U171 ( .A(n191), .Z(n186) );
  GTECH_NOT U172 ( .A(n175), .Z(n185) );
  GTECH_NAND2 U173 ( .A(I_b[7]), .B(I_a[3]), .Z(n175) );
  GTECH_NOT U174 ( .A(n173), .Z(n176) );
  GTECH_NAND2 U175 ( .A(I_b[6]), .B(I_a[4]), .Z(n173) );
  GTECH_OAI22 U176 ( .A(n192), .B(n193), .C(n194), .D(n195), .Z(n181) );
  GTECH_AND_NOT U177 ( .A(n192), .B(n196), .Z(n194) );
  GTECH_NOT U178 ( .A(n180), .Z(n169) );
  GTECH_NAND2 U179 ( .A(I_a[5]), .B(I_b[5]), .Z(n180) );
  GTECH_ADD_ABC U180 ( .A(n197), .B(n198), .C(n199), .COUT(n164) );
  GTECH_NOT U181 ( .A(n200), .Z(n199) );
  GTECH_XOR3 U182 ( .A(n196), .B(n201), .C(n192), .Z(n198) );
  GTECH_NOT U183 ( .A(n202), .Z(n192) );
  GTECH_NOT U184 ( .A(n157), .Z(n183) );
  GTECH_XOR2 U185 ( .A(n182), .B(n154), .Z(n157) );
  GTECH_AOI2N2 U186 ( .A(n203), .B(n204), .C(n205), .D(n206), .Z(n154) );
  GTECH_NAND2 U187 ( .A(n205), .B(n206), .Z(n204) );
  GTECH_XOR2 U188 ( .A(n207), .B(n152), .Z(n182) );
  GTECH_OA21 U189 ( .A(n208), .B(n209), .C(n210), .Z(n152) );
  GTECH_AO21 U190 ( .A(n208), .B(n209), .C(n211), .Z(n210) );
  GTECH_NOT U191 ( .A(n212), .Z(n208) );
  GTECH_NAND2 U192 ( .A(I_a[7]), .B(I_b[3]), .Z(n207) );
  GTECH_OA21 U193 ( .A(n213), .B(n214), .C(n215), .Z(n156) );
  GTECH_AO21 U194 ( .A(n213), .B(n214), .C(n216), .Z(n215) );
  GTECH_XOR3 U195 ( .A(n213), .B(n217), .C(n216), .Z(N149) );
  GTECH_XOR2 U196 ( .A(n197), .B(n218), .Z(n216) );
  GTECH_XOR4 U197 ( .A(n201), .B(n202), .C(n200), .D(n196), .Z(n218) );
  GTECH_NOT U198 ( .A(n193), .Z(n196) );
  GTECH_NAND2 U199 ( .A(I_a[5]), .B(I_b[4]), .Z(n193) );
  GTECH_XOR3 U200 ( .A(n190), .B(n219), .C(n191), .Z(n200) );
  GTECH_AO21 U201 ( .A(n220), .B(n221), .C(n222), .Z(n191) );
  GTECH_NOT U202 ( .A(n223), .Z(n222) );
  GTECH_NOT U203 ( .A(n189), .Z(n219) );
  GTECH_NAND2 U204 ( .A(I_b[7]), .B(I_a[2]), .Z(n189) );
  GTECH_NOT U205 ( .A(n187), .Z(n190) );
  GTECH_NAND2 U206 ( .A(I_b[6]), .B(I_a[3]), .Z(n187) );
  GTECH_OAI22 U207 ( .A(n224), .B(n225), .C(n226), .D(n227), .Z(n202) );
  GTECH_AND_NOT U208 ( .A(n224), .B(n228), .Z(n226) );
  GTECH_NOT U209 ( .A(n195), .Z(n201) );
  GTECH_NAND2 U210 ( .A(I_b[5]), .B(I_a[4]), .Z(n195) );
  GTECH_ADD_ABC U211 ( .A(n229), .B(n230), .C(n231), .COUT(n197) );
  GTECH_XOR3 U212 ( .A(n228), .B(n232), .C(n224), .Z(n230) );
  GTECH_NOT U213 ( .A(n233), .Z(n224) );
  GTECH_NOT U214 ( .A(n225), .Z(n228) );
  GTECH_OA21 U215 ( .A(n234), .B(n235), .C(n236), .Z(n229) );
  GTECH_AO21 U216 ( .A(n234), .B(n235), .C(n237), .Z(n236) );
  GTECH_NOT U217 ( .A(n214), .Z(n217) );
  GTECH_XOR3 U218 ( .A(n238), .B(n205), .C(n203), .Z(n214) );
  GTECH_XOR3 U219 ( .A(n239), .B(n240), .C(n212), .Z(n203) );
  GTECH_OAI22 U220 ( .A(n241), .B(n242), .C(n243), .D(n244), .Z(n212) );
  GTECH_AND_NOT U221 ( .A(n241), .B(n245), .Z(n243) );
  GTECH_NOT U222 ( .A(n246), .Z(n241) );
  GTECH_NOT U223 ( .A(n211), .Z(n240) );
  GTECH_NAND2 U224 ( .A(I_a[6]), .B(I_b[3]), .Z(n211) );
  GTECH_NOT U225 ( .A(n209), .Z(n239) );
  GTECH_NAND2 U226 ( .A(I_a[7]), .B(I_b[2]), .Z(n209) );
  GTECH_ADD_ABC U227 ( .A(n247), .B(n248), .C(n249), .COUT(n205) );
  GTECH_XOR2 U228 ( .A(n250), .B(n251), .Z(n248) );
  GTECH_AND_NOT U229 ( .A(I_a[7]), .B(n252), .Z(n251) );
  GTECH_NOT U230 ( .A(I_b[1]), .Z(n252) );
  GTECH_NOT U231 ( .A(n253), .Z(n250) );
  GTECH_NOT U232 ( .A(n206), .Z(n238) );
  GTECH_NAND2 U233 ( .A(I_a[7]), .B(n253), .Z(n206) );
  GTECH_ADD_ABC U234 ( .A(n254), .B(n255), .C(n256), .COUT(n213) );
  GTECH_XOR3 U235 ( .A(n247), .B(n257), .C(n249), .Z(n255) );
  GTECH_NOT U236 ( .A(n258), .Z(n249) );
  GTECH_XOR2 U237 ( .A(n254), .B(n259), .Z(N148) );
  GTECH_XOR4 U238 ( .A(n257), .B(n258), .C(n256), .D(n247), .Z(n259) );
  GTECH_ADD_ABC U239 ( .A(n260), .B(n261), .C(n262), .COUT(n247) );
  GTECH_XOR3 U240 ( .A(n263), .B(n264), .C(n265), .Z(n261) );
  GTECH_XOR2 U241 ( .A(n266), .B(n267), .Z(n256) );
  GTECH_OA22 U242 ( .A(n268), .B(n237), .C(n234), .D(n235), .Z(n267) );
  GTECH_AND_NOT U243 ( .A(n234), .B(n269), .Z(n268) );
  GTECH_XOR4 U244 ( .A(n232), .B(n233), .C(n225), .D(n231), .Z(n266) );
  GTECH_XOR3 U245 ( .A(n221), .B(n220), .C(n223), .Z(n231) );
  GTECH_NAND3 U246 ( .A(I_b[6]), .B(I_a[1]), .C(n270), .Z(n223) );
  GTECH_NOT U247 ( .A(n271), .Z(n220) );
  GTECH_NAND2 U248 ( .A(I_b[7]), .B(I_a[1]), .Z(n271) );
  GTECH_NOT U249 ( .A(n272), .Z(n221) );
  GTECH_NAND2 U250 ( .A(I_b[6]), .B(I_a[2]), .Z(n272) );
  GTECH_NAND2 U251 ( .A(I_b[4]), .B(I_a[4]), .Z(n225) );
  GTECH_OAI22 U252 ( .A(n273), .B(n274), .C(n275), .D(n276), .Z(n233) );
  GTECH_AND_NOT U253 ( .A(n273), .B(n277), .Z(n275) );
  GTECH_NOT U254 ( .A(n278), .Z(n273) );
  GTECH_NOT U255 ( .A(n227), .Z(n232) );
  GTECH_NAND2 U256 ( .A(I_b[5]), .B(I_a[3]), .Z(n227) );
  GTECH_XOR3 U257 ( .A(n245), .B(n279), .C(n246), .Z(n258) );
  GTECH_OAI22 U258 ( .A(n280), .B(n281), .C(n282), .D(n283), .Z(n246) );
  GTECH_AND_NOT U259 ( .A(n280), .B(n284), .Z(n282) );
  GTECH_NOT U260 ( .A(n285), .Z(n280) );
  GTECH_NOT U261 ( .A(n244), .Z(n279) );
  GTECH_NAND2 U262 ( .A(I_a[5]), .B(I_b[3]), .Z(n244) );
  GTECH_NOT U263 ( .A(n242), .Z(n245) );
  GTECH_NAND2 U264 ( .A(I_a[6]), .B(I_b[2]), .Z(n242) );
  GTECH_XOR2 U265 ( .A(n286), .B(n253), .Z(n257) );
  GTECH_OAI22 U266 ( .A(n265), .B(n287), .C(n288), .D(n289), .Z(n253) );
  GTECH_AND_NOT U267 ( .A(n265), .B(n263), .Z(n288) );
  GTECH_NOT U268 ( .A(n290), .Z(n265) );
  GTECH_NAND2 U269 ( .A(I_a[7]), .B(I_b[1]), .Z(n286) );
  GTECH_ADD_ABC U270 ( .A(n291), .B(n292), .C(n293), .COUT(n254) );
  GTECH_NOT U271 ( .A(n294), .Z(n293) );
  GTECH_XOR3 U272 ( .A(n260), .B(n295), .C(n262), .Z(n292) );
  GTECH_NOT U273 ( .A(n296), .Z(n262) );
  GTECH_NOT U274 ( .A(n297), .Z(n295) );
  GTECH_XOR2 U275 ( .A(n298), .B(n291), .Z(N147) );
  GTECH_ADD_ABC U276 ( .A(n299), .B(n300), .C(n301), .COUT(n291) );
  GTECH_XOR3 U277 ( .A(n302), .B(n303), .C(n304), .Z(n300) );
  GTECH_OA21 U278 ( .A(n305), .B(n306), .C(n307), .Z(n299) );
  GTECH_AO21 U279 ( .A(n305), .B(n306), .C(n308), .Z(n307) );
  GTECH_XOR4 U280 ( .A(n296), .B(n260), .C(n297), .D(n294), .Z(n298) );
  GTECH_XOR3 U281 ( .A(n309), .B(n235), .C(n234), .Z(n294) );
  GTECH_XOR2 U282 ( .A(n310), .B(n270), .Z(n234) );
  GTECH_NOT U283 ( .A(n311), .Z(n270) );
  GTECH_NAND2 U284 ( .A(I_b[7]), .B(I_a[0]), .Z(n311) );
  GTECH_NAND2 U285 ( .A(I_b[6]), .B(I_a[1]), .Z(n310) );
  GTECH_NOT U286 ( .A(n269), .Z(n235) );
  GTECH_XOR3 U287 ( .A(n277), .B(n312), .C(n278), .Z(n269) );
  GTECH_AO21 U288 ( .A(n313), .B(n314), .C(n315), .Z(n278) );
  GTECH_NOT U289 ( .A(n316), .Z(n315) );
  GTECH_NOT U290 ( .A(n276), .Z(n312) );
  GTECH_NAND2 U291 ( .A(I_b[5]), .B(I_a[2]), .Z(n276) );
  GTECH_NOT U292 ( .A(n274), .Z(n277) );
  GTECH_NAND2 U293 ( .A(I_b[4]), .B(I_a[3]), .Z(n274) );
  GTECH_NOT U294 ( .A(n237), .Z(n309) );
  GTECH_NAND3 U295 ( .A(I_a[0]), .B(n317), .C(I_b[6]), .Z(n237) );
  GTECH_NOT U296 ( .A(n318), .Z(n317) );
  GTECH_XOR3 U297 ( .A(n263), .B(n264), .C(n290), .Z(n297) );
  GTECH_OAI22 U298 ( .A(n319), .B(n320), .C(n321), .D(n322), .Z(n290) );
  GTECH_AND_NOT U299 ( .A(n319), .B(n323), .Z(n321) );
  GTECH_NOT U300 ( .A(n289), .Z(n264) );
  GTECH_NAND2 U301 ( .A(I_a[6]), .B(I_b[1]), .Z(n289) );
  GTECH_NOT U302 ( .A(n287), .Z(n263) );
  GTECH_NAND2 U303 ( .A(I_a[7]), .B(I_b[0]), .Z(n287) );
  GTECH_ADD_ABC U304 ( .A(n302), .B(n324), .C(n304), .COUT(n260) );
  GTECH_NOT U305 ( .A(n325), .Z(n304) );
  GTECH_XOR3 U306 ( .A(n323), .B(n326), .C(n319), .Z(n324) );
  GTECH_NOT U307 ( .A(n327), .Z(n319) );
  GTECH_XOR3 U308 ( .A(n284), .B(n328), .C(n285), .Z(n296) );
  GTECH_OAI22 U309 ( .A(n329), .B(n330), .C(n331), .D(n332), .Z(n285) );
  GTECH_AND_NOT U310 ( .A(n329), .B(n333), .Z(n331) );
  GTECH_NOT U311 ( .A(n334), .Z(n329) );
  GTECH_NOT U312 ( .A(n283), .Z(n328) );
  GTECH_NAND2 U313 ( .A(I_b[3]), .B(I_a[4]), .Z(n283) );
  GTECH_NOT U314 ( .A(n281), .Z(n284) );
  GTECH_NAND2 U315 ( .A(I_a[5]), .B(I_b[2]), .Z(n281) );
  GTECH_XOR2 U316 ( .A(n335), .B(n336), .Z(N146) );
  GTECH_XOR4 U317 ( .A(n303), .B(n325), .C(n301), .D(n302), .Z(n336) );
  GTECH_ADD_ABC U318 ( .A(n337), .B(n338), .C(n339), .COUT(n302) );
  GTECH_NOT U319 ( .A(n340), .Z(n339) );
  GTECH_XOR3 U320 ( .A(n341), .B(n342), .C(n343), .Z(n338) );
  GTECH_XOR2 U321 ( .A(n318), .B(n344), .Z(n301) );
  GTECH_AND_NOT U322 ( .A(I_b[6]), .B(n345), .Z(n344) );
  GTECH_XOR3 U323 ( .A(n314), .B(n313), .C(n316), .Z(n318) );
  GTECH_NAND3 U324 ( .A(I_b[4]), .B(I_a[1]), .C(n346), .Z(n316) );
  GTECH_NOT U325 ( .A(n347), .Z(n313) );
  GTECH_NAND2 U326 ( .A(I_b[5]), .B(I_a[1]), .Z(n347) );
  GTECH_NOT U327 ( .A(n348), .Z(n314) );
  GTECH_NAND2 U328 ( .A(I_b[4]), .B(I_a[2]), .Z(n348) );
  GTECH_XOR3 U329 ( .A(n333), .B(n349), .C(n334), .Z(n325) );
  GTECH_OAI22 U330 ( .A(n350), .B(n351), .C(n352), .D(n353), .Z(n334) );
  GTECH_AND_NOT U331 ( .A(n350), .B(n354), .Z(n352) );
  GTECH_NOT U332 ( .A(n355), .Z(n350) );
  GTECH_NOT U333 ( .A(n332), .Z(n349) );
  GTECH_NAND2 U334 ( .A(I_b[3]), .B(I_a[3]), .Z(n332) );
  GTECH_NOT U335 ( .A(n330), .Z(n333) );
  GTECH_NAND2 U336 ( .A(I_b[2]), .B(I_a[4]), .Z(n330) );
  GTECH_NOT U337 ( .A(n356), .Z(n303) );
  GTECH_XOR3 U338 ( .A(n323), .B(n326), .C(n327), .Z(n356) );
  GTECH_OAI22 U339 ( .A(n343), .B(n357), .C(n358), .D(n359), .Z(n327) );
  GTECH_AND_NOT U340 ( .A(n343), .B(n341), .Z(n358) );
  GTECH_NOT U341 ( .A(n357), .Z(n341) );
  GTECH_NOT U342 ( .A(n360), .Z(n343) );
  GTECH_NOT U343 ( .A(n322), .Z(n326) );
  GTECH_NAND2 U344 ( .A(I_a[5]), .B(I_b[1]), .Z(n322) );
  GTECH_NOT U345 ( .A(n320), .Z(n323) );
  GTECH_NAND2 U346 ( .A(I_a[6]), .B(I_b[0]), .Z(n320) );
  GTECH_OA22 U347 ( .A(n361), .B(n308), .C(n305), .D(n306), .Z(n335) );
  GTECH_AND_NOT U348 ( .A(n305), .B(n362), .Z(n361) );
  GTECH_XOR3 U349 ( .A(n363), .B(n306), .C(n305), .Z(N145) );
  GTECH_XOR2 U350 ( .A(n364), .B(n346), .Z(n305) );
  GTECH_NOT U351 ( .A(n365), .Z(n346) );
  GTECH_NAND2 U352 ( .A(I_b[5]), .B(I_a[0]), .Z(n365) );
  GTECH_NAND2 U353 ( .A(I_b[4]), .B(I_a[1]), .Z(n364) );
  GTECH_NOT U354 ( .A(n362), .Z(n306) );
  GTECH_XOR2 U355 ( .A(n366), .B(n337), .Z(n362) );
  GTECH_ADD_ABC U356 ( .A(n367), .B(n368), .C(n369), .COUT(n337) );
  GTECH_XOR3 U357 ( .A(n370), .B(n371), .C(n372), .Z(n368) );
  GTECH_OA21 U358 ( .A(n373), .B(n374), .C(n375), .Z(n367) );
  GTECH_AO21 U359 ( .A(n373), .B(n374), .C(n376), .Z(n375) );
  GTECH_XOR4 U360 ( .A(n342), .B(n360), .C(n357), .D(n340), .Z(n366) );
  GTECH_XOR3 U361 ( .A(n354), .B(n377), .C(n355), .Z(n340) );
  GTECH_AO21 U362 ( .A(n378), .B(n379), .C(n380), .Z(n355) );
  GTECH_NOT U363 ( .A(n381), .Z(n380) );
  GTECH_NOT U364 ( .A(n353), .Z(n377) );
  GTECH_NAND2 U365 ( .A(I_b[3]), .B(I_a[2]), .Z(n353) );
  GTECH_NOT U366 ( .A(n351), .Z(n354) );
  GTECH_NAND2 U367 ( .A(I_b[2]), .B(I_a[3]), .Z(n351) );
  GTECH_NAND2 U368 ( .A(I_a[5]), .B(I_b[0]), .Z(n357) );
  GTECH_OAI22 U369 ( .A(n372), .B(n382), .C(n383), .D(n384), .Z(n360) );
  GTECH_AND_NOT U370 ( .A(n372), .B(n370), .Z(n383) );
  GTECH_NOT U371 ( .A(n385), .Z(n372) );
  GTECH_NOT U372 ( .A(n359), .Z(n342) );
  GTECH_NAND2 U373 ( .A(I_a[4]), .B(I_b[1]), .Z(n359) );
  GTECH_NOT U374 ( .A(n308), .Z(n363) );
  GTECH_NAND3 U375 ( .A(I_a[0]), .B(n386), .C(I_b[4]), .Z(n308) );
  GTECH_XOR2 U376 ( .A(n387), .B(n386), .Z(N144) );
  GTECH_XOR2 U377 ( .A(n388), .B(n389), .Z(n386) );
  GTECH_XOR4 U378 ( .A(n371), .B(n385), .C(n369), .D(n370), .Z(n389) );
  GTECH_NOT U379 ( .A(n382), .Z(n370) );
  GTECH_NAND2 U380 ( .A(I_a[4]), .B(I_b[0]), .Z(n382) );
  GTECH_XOR3 U381 ( .A(n379), .B(n378), .C(n381), .Z(n369) );
  GTECH_NAND3 U382 ( .A(I_b[2]), .B(I_a[1]), .C(n390), .Z(n381) );
  GTECH_NOT U383 ( .A(n391), .Z(n378) );
  GTECH_NAND2 U384 ( .A(I_b[3]), .B(I_a[1]), .Z(n391) );
  GTECH_NOT U385 ( .A(n392), .Z(n379) );
  GTECH_NAND2 U386 ( .A(I_b[2]), .B(I_a[2]), .Z(n392) );
  GTECH_OAI22 U387 ( .A(n393), .B(n394), .C(n395), .D(n396), .Z(n385) );
  GTECH_AND_NOT U388 ( .A(n393), .B(n397), .Z(n395) );
  GTECH_NOT U389 ( .A(n398), .Z(n393) );
  GTECH_NOT U390 ( .A(n384), .Z(n371) );
  GTECH_NAND2 U391 ( .A(I_a[3]), .B(I_b[1]), .Z(n384) );
  GTECH_OA22 U392 ( .A(n399), .B(n376), .C(n373), .D(n374), .Z(n388) );
  GTECH_AND_NOT U393 ( .A(n373), .B(n400), .Z(n399) );
  GTECH_AND_NOT U394 ( .A(I_b[4]), .B(n345), .Z(n387) );
  GTECH_XOR3 U395 ( .A(n401), .B(n374), .C(n373), .Z(N143) );
  GTECH_XOR2 U396 ( .A(n402), .B(n390), .Z(n373) );
  GTECH_NOT U397 ( .A(n403), .Z(n390) );
  GTECH_NAND2 U398 ( .A(I_b[3]), .B(I_a[0]), .Z(n403) );
  GTECH_NAND2 U399 ( .A(I_b[2]), .B(I_a[1]), .Z(n402) );
  GTECH_NOT U400 ( .A(n400), .Z(n374) );
  GTECH_XOR3 U401 ( .A(n397), .B(n404), .C(n398), .Z(n400) );
  GTECH_AO21 U402 ( .A(n405), .B(n406), .C(n407), .Z(n398) );
  GTECH_NOT U403 ( .A(n408), .Z(n407) );
  GTECH_NOT U404 ( .A(n396), .Z(n404) );
  GTECH_NAND2 U405 ( .A(I_b[1]), .B(I_a[2]), .Z(n396) );
  GTECH_NOT U406 ( .A(n394), .Z(n397) );
  GTECH_NAND2 U407 ( .A(I_b[0]), .B(I_a[3]), .Z(n394) );
  GTECH_NOT U408 ( .A(n376), .Z(n401) );
  GTECH_NAND3 U409 ( .A(I_a[0]), .B(n409), .C(I_b[2]), .Z(n376) );
  GTECH_XOR2 U410 ( .A(n410), .B(n409), .Z(N142) );
  GTECH_NOT U411 ( .A(n411), .Z(n409) );
  GTECH_XOR3 U412 ( .A(n405), .B(n406), .C(n408), .Z(n411) );
  GTECH_NAND3 U413 ( .A(n412), .B(I_b[0]), .C(I_a[1]), .Z(n408) );
  GTECH_NOT U414 ( .A(n413), .Z(n406) );
  GTECH_NAND2 U415 ( .A(I_a[1]), .B(I_b[1]), .Z(n413) );
  GTECH_NOT U416 ( .A(n414), .Z(n405) );
  GTECH_NAND2 U417 ( .A(I_b[0]), .B(I_a[2]), .Z(n414) );
  GTECH_AND_NOT U418 ( .A(I_b[2]), .B(n345), .Z(n410) );
  GTECH_NOT U419 ( .A(I_a[0]), .Z(n345) );
  GTECH_XOR2 U420 ( .A(n412), .B(n415), .Z(N141) );
  GTECH_AND_NOT U421 ( .A(I_a[1]), .B(n416), .Z(n415) );
  GTECH_NOT U422 ( .A(n417), .Z(n412) );
  GTECH_NAND2 U423 ( .A(I_a[0]), .B(I_b[1]), .Z(n417) );
  GTECH_AND_NOT U424 ( .A(I_a[0]), .B(n416), .Z(N140) );
  GTECH_NOT U425 ( .A(I_b[0]), .Z(n416) );
endmodule

