
module fraction_multiplier4 ( CLK, St, Mplier, Mcand, Product, Done );
  input [3:0] Mplier;
  input [3:0] Mcand;
  output [6:0] Product;
  input CLK, St;
  output Done;
  wire   N40, N41, N42, N44, N46, N48, N50, N52, N54, N56, N57, N58, N63, n12,
         n14, n15, n16, n17, n18, n19, n76, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143;
  wire   [2:0] State;

  GTECH_FD1 State_reg_0_ ( .D(N40), .CP(CLK), .Q(State[0]), .QN(n86) );
  GTECH_FD1 State_reg_1_ ( .D(N41), .CP(CLK), .Q(State[1]), .QN(n85) );
  GTECH_FD1 State_reg_2_ ( .D(N42), .CP(CLK), .Q(State[2]), .QN(n87) );
  GTECH_FJK1S B_reg_0_ ( .J(n76), .K(n76), .TI(N52), .TE(N57), .CP(CLK), .Q(
        Product[0]), .QN(n12) );
  GTECH_FJK1S A_reg_3_ ( .J(n76), .K(n76), .TI(N50), .TE(N63), .CP(CLK), .QN(
        n84) );
  GTECH_FJK1S A_reg_0_ ( .J(n76), .K(n76), .TI(N44), .TE(N57), .CP(CLK), .Q(
        Product[4]), .QN(n14) );
  GTECH_FJK1S A_reg_1_ ( .J(n76), .K(n76), .TI(N46), .TE(N57), .CP(CLK), .Q(
        Product[5]), .QN(n15) );
  GTECH_FJK1S A_reg_2_ ( .J(n76), .K(n76), .TI(N48), .TE(N57), .CP(CLK), .Q(
        Product[6]), .QN(n16) );
  GTECH_FJK1S B_reg_3_ ( .J(n76), .K(n76), .TI(N58), .TE(N57), .CP(CLK), .Q(
        Product[3]), .QN(n17) );
  GTECH_FJK1S B_reg_2_ ( .J(n76), .K(n76), .TI(N56), .TE(N57), .CP(CLK), .Q(
        Product[2]), .QN(n18) );
  GTECH_FJK1S B_reg_1_ ( .J(n76), .K(n76), .TI(N54), .TE(N57), .CP(CLK), .Q(
        Product[1]), .QN(n19) );
  GTECH_ZERO U81 ( .Z(n76) );
  GTECH_AND2 U82 ( .A(N57), .B(n88), .Z(N63) );
  GTECH_NOT U83 ( .A(n89), .Z(N58) );
  GTECH_AOI222 U84 ( .A(Mplier[3]), .B(n90), .C(n91), .D(n92), .E(n93), .F(n94), .Z(n89) );
  GTECH_NOT U85 ( .A(n14), .Z(n94) );
  GTECH_OAI21 U86 ( .A(Mcand[0]), .B(n95), .C(n88), .Z(n93) );
  GTECH_AND_NOT U87 ( .A(n96), .B(n12), .Z(n91) );
  GTECH_AO21 U88 ( .A(n90), .B(St), .C(n96), .Z(N57) );
  GTECH_NOT U89 ( .A(n95), .Z(n96) );
  GTECH_OAI2N2 U90 ( .A(n17), .B(n95), .C(Mplier[2]), .D(n90), .Z(N56) );
  GTECH_OAI2N2 U91 ( .A(n18), .B(n95), .C(Mplier[1]), .D(n90), .Z(N54) );
  GTECH_OAI2N2 U92 ( .A(n19), .B(n95), .C(Mplier[0]), .D(n90), .Z(N52) );
  GTECH_MUX2 U93 ( .A(n97), .B(n98), .S(Mcand[3]), .Z(N50) );
  GTECH_MUX2 U94 ( .A(n99), .B(n100), .S(n84), .Z(N48) );
  GTECH_MUX2 U95 ( .A(n101), .B(n102), .S(Mcand[3]), .Z(n100) );
  GTECH_OR_NOT U96 ( .A(n103), .B(n88), .Z(n99) );
  GTECH_MUX2 U97 ( .A(n102), .B(n101), .S(Mcand[3]), .Z(n103) );
  GTECH_OAI22 U98 ( .A(n104), .B(n105), .C(n106), .D(n107), .Z(n101) );
  GTECH_AO22 U99 ( .A(n105), .B(n108), .C(n107), .D(n109), .Z(n102) );
  GTECH_OAI21 U100 ( .A(Mcand[2]), .B(n110), .C(n111), .Z(n107) );
  GTECH_AO21 U101 ( .A(n110), .B(Mcand[2]), .C(n112), .Z(n111) );
  GTECH_OAI21 U102 ( .A(Mcand[2]), .B(n113), .C(n114), .Z(n105) );
  GTECH_AO21 U103 ( .A(n113), .B(Mcand[2]), .C(n16), .Z(n114) );
  GTECH_MUX2 U104 ( .A(n115), .B(n116), .S(n112), .Z(N46) );
  GTECH_NOT U105 ( .A(n16), .Z(n112) );
  GTECH_NAND2 U106 ( .A(n117), .B(n88), .Z(n116) );
  GTECH_MUX2 U107 ( .A(n118), .B(n119), .S(Mcand[2]), .Z(n117) );
  GTECH_NOT U108 ( .A(n120), .Z(n115) );
  GTECH_MUX2 U109 ( .A(n119), .B(n118), .S(Mcand[2]), .Z(n120) );
  GTECH_AOI2N2 U110 ( .A(n121), .B(n109), .C(n113), .D(n104), .Z(n118) );
  GTECH_NOT U111 ( .A(n122), .Z(n113) );
  GTECH_NOT U112 ( .A(n110), .Z(n121) );
  GTECH_AOI2N2 U113 ( .A(n110), .B(n109), .C(n122), .D(n104), .Z(n119) );
  GTECH_ADD_ABC U114 ( .A(n123), .B(n124), .C(n125), .COUT(n122) );
  GTECH_NAND2 U115 ( .A(Mcand[0]), .B(n14), .Z(n123) );
  GTECH_OAI21 U116 ( .A(n15), .B(n124), .C(n126), .Z(n110) );
  GTECH_OR3 U117 ( .A(n127), .B(n14), .C(n128), .Z(n126) );
  GTECH_AO21 U118 ( .A(n129), .B(n127), .C(n130), .Z(N44) );
  GTECH_NOT U119 ( .A(n131), .Z(n130) );
  GTECH_MUX2 U120 ( .A(n132), .B(n133), .S(n15), .Z(n131) );
  GTECH_NAND2 U121 ( .A(Mcand[1]), .B(n134), .Z(n133) );
  GTECH_AND_NOT U122 ( .A(n88), .B(n135), .Z(n132) );
  GTECH_MUX2 U123 ( .A(n134), .B(n129), .S(Mcand[1]), .Z(n135) );
  GTECH_OAI21 U124 ( .A(n92), .B(n104), .C(n136), .Z(n134) );
  GTECH_OAI21 U125 ( .A(n14), .B(n128), .C(n109), .Z(n136) );
  GTECH_NOT U126 ( .A(n108), .Z(n104) );
  GTECH_OR_NOT U127 ( .A(n95), .B(n12), .Z(n88) );
  GTECH_AND_NOT U128 ( .A(n137), .B(n97), .Z(n95) );
  GTECH_AND_NOT U129 ( .A(n124), .B(n125), .Z(n127) );
  GTECH_NOT U130 ( .A(n15), .Z(n125) );
  GTECH_NOT U131 ( .A(Mcand[1]), .Z(n124) );
  GTECH_AO21 U132 ( .A(n92), .B(n108), .C(n138), .Z(n129) );
  GTECH_NOR3 U133 ( .A(n128), .B(n14), .C(n106), .Z(n138) );
  GTECH_NOT U134 ( .A(n109), .Z(n106) );
  GTECH_AND_NOT U135 ( .A(n98), .B(n12), .Z(n109) );
  GTECH_AND_NOT U136 ( .A(n97), .B(n12), .Z(n108) );
  GTECH_AND_NOT U137 ( .A(n14), .B(n128), .Z(n92) );
  GTECH_NOT U138 ( .A(Mcand[0]), .Z(n128) );
  GTECH_OR_NOT U139 ( .A(n97), .B(n139), .Z(N42) );
  GTECH_NAND3 U140 ( .A(n140), .B(n141), .C(n98), .Z(n139) );
  GTECH_AOI21 U141 ( .A(n141), .B(n140), .C(n137), .Z(N41) );
  GTECH_NOT U142 ( .A(n98), .Z(n137) );
  GTECH_NOT U143 ( .A(n86), .Z(n141) );
  GTECH_AO21 U144 ( .A(n90), .B(St), .C(n142), .Z(N40) );
  GTECH_AO21 U145 ( .A(n98), .B(n86), .C(n97), .Z(n142) );
  GTECH_AND_NOT U146 ( .A(n143), .B(n87), .Z(n97) );
  GTECH_AND_NOT U147 ( .A(n87), .B(n143), .Z(n98) );
  GTECH_AND2 U148 ( .A(n87), .B(n143), .Z(n90) );
  GTECH_AND2 U149 ( .A(n86), .B(n85), .Z(n143) );
  GTECH_NOR3 U150 ( .A(n86), .B(n87), .C(n140), .Z(Done) );
  GTECH_NOT U151 ( .A(n85), .Z(n140) );
endmodule

