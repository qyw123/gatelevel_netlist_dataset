
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370;

  GTECH_MUX2 U123 ( .A(n262), .B(n263), .S(n264), .Z(sum[9]) );
  GTECH_OA21 U124 ( .A(n265), .B(n266), .C(n267), .Z(n264) );
  GTECH_OAI21 U125 ( .A(a[8]), .B(n268), .C(b[8]), .Z(n267) );
  GTECH_XOR2 U126 ( .A(b[9]), .B(a[9]), .Z(n263) );
  GTECH_NAND2 U127 ( .A(n269), .B(n270), .Z(n262) );
  GTECH_XOR2 U128 ( .A(n268), .B(n271), .Z(sum[8]) );
  GTECH_MUX2 U129 ( .A(n272), .B(n273), .S(n274), .Z(sum[7]) );
  GTECH_XNOR2 U130 ( .A(n275), .B(n276), .Z(n273) );
  GTECH_XOR2 U131 ( .A(n275), .B(n277), .Z(n272) );
  GTECH_OA21 U132 ( .A(n278), .B(n279), .C(n280), .Z(n277) );
  GTECH_NOT U133 ( .A(n281), .Z(n279) );
  GTECH_XNOR2 U134 ( .A(a[7]), .B(b[7]), .Z(n275) );
  GTECH_MUX2 U135 ( .A(n282), .B(n283), .S(n274), .Z(sum[6]) );
  GTECH_XNOR2 U136 ( .A(n284), .B(n285), .Z(n283) );
  GTECH_XOR2 U137 ( .A(n284), .B(n281), .Z(n282) );
  GTECH_AO21 U138 ( .A(n286), .B(n287), .C(n288), .Z(n281) );
  GTECH_AND_NOT U139 ( .A(n280), .B(n278), .Z(n284) );
  GTECH_MUX2 U140 ( .A(n289), .B(n290), .S(n291), .Z(sum[5]) );
  GTECH_AND_NOT U141 ( .A(n286), .B(n288), .Z(n291) );
  GTECH_OAI21 U142 ( .A(n287), .B(n274), .C(n292), .Z(n290) );
  GTECH_AO21 U143 ( .A(n292), .B(n274), .C(n287), .Z(n289) );
  GTECH_XOR2 U144 ( .A(n274), .B(n293), .Z(sum[4]) );
  GTECH_MUX2 U145 ( .A(n294), .B(n295), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U146 ( .A(n296), .B(n297), .Z(n295) );
  GTECH_XOR2 U147 ( .A(n296), .B(n298), .Z(n294) );
  GTECH_AO21 U148 ( .A(n299), .B(n300), .C(n301), .Z(n298) );
  GTECH_XOR2 U149 ( .A(a[3]), .B(b[3]), .Z(n296) );
  GTECH_MUX2 U150 ( .A(n302), .B(n303), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U151 ( .A(n304), .B(n305), .Z(n303) );
  GTECH_XOR2 U152 ( .A(n304), .B(n300), .Z(n302) );
  GTECH_AO21 U153 ( .A(n306), .B(n307), .C(n308), .Z(n300) );
  GTECH_AND_NOT U154 ( .A(n299), .B(n301), .Z(n304) );
  GTECH_MUX2 U155 ( .A(n309), .B(n310), .S(n311), .Z(sum[1]) );
  GTECH_AND_NOT U156 ( .A(n306), .B(n308), .Z(n311) );
  GTECH_OAI21 U157 ( .A(cin), .B(n307), .C(n312), .Z(n310) );
  GTECH_AO21 U158 ( .A(n312), .B(cin), .C(n307), .Z(n309) );
  GTECH_MUX2 U159 ( .A(n313), .B(n314), .S(n315), .Z(sum[15]) );
  GTECH_XOR2 U160 ( .A(n316), .B(n317), .Z(n314) );
  GTECH_XOR2 U161 ( .A(n316), .B(n318), .Z(n313) );
  GTECH_AND2 U162 ( .A(n319), .B(n320), .Z(n318) );
  GTECH_AO21 U163 ( .A(n321), .B(n322), .C(n323), .Z(n319) );
  GTECH_XNOR2 U164 ( .A(a[15]), .B(b[15]), .Z(n316) );
  GTECH_MUX2 U165 ( .A(n324), .B(n325), .S(n315), .Z(sum[14]) );
  GTECH_XNOR2 U166 ( .A(n326), .B(n327), .Z(n325) );
  GTECH_XNOR2 U167 ( .A(n326), .B(n323), .Z(n324) );
  GTECH_AOI22 U168 ( .A(a[13]), .B(b[13]), .C(n328), .D(n329), .Z(n323) );
  GTECH_NOT U169 ( .A(n330), .Z(n328) );
  GTECH_OA21 U170 ( .A(b[14]), .B(a[14]), .C(n320), .Z(n326) );
  GTECH_MUX2 U171 ( .A(n331), .B(n332), .S(n315), .Z(sum[13]) );
  GTECH_XOR2 U172 ( .A(n333), .B(n334), .Z(n332) );
  GTECH_XNOR2 U173 ( .A(n329), .B(n334), .Z(n331) );
  GTECH_AO21 U174 ( .A(a[13]), .B(b[13]), .C(n330), .Z(n334) );
  GTECH_NAND2 U175 ( .A(n335), .B(n336), .Z(sum[12]) );
  GTECH_OAI21 U176 ( .A(n329), .B(n333), .C(n315), .Z(n335) );
  GTECH_MUX2 U177 ( .A(n337), .B(n338), .S(n265), .Z(sum[11]) );
  GTECH_XNOR2 U178 ( .A(n339), .B(n340), .Z(n338) );
  GTECH_AND2 U179 ( .A(n341), .B(n342), .Z(n340) );
  GTECH_AO21 U180 ( .A(n343), .B(n344), .C(n345), .Z(n341) );
  GTECH_XOR2 U181 ( .A(n339), .B(n346), .Z(n337) );
  GTECH_XOR2 U182 ( .A(a[11]), .B(b[11]), .Z(n339) );
  GTECH_MUX2 U183 ( .A(n347), .B(n348), .S(n265), .Z(sum[10]) );
  GTECH_XNOR2 U184 ( .A(n349), .B(n345), .Z(n348) );
  GTECH_AND2 U185 ( .A(n350), .B(n269), .Z(n345) );
  GTECH_NOT U186 ( .A(n351), .Z(n269) );
  GTECH_NAND3 U187 ( .A(b[8]), .B(n270), .C(a[8]), .Z(n350) );
  GTECH_XNOR2 U188 ( .A(n349), .B(n352), .Z(n347) );
  GTECH_OA21 U189 ( .A(b[10]), .B(a[10]), .C(n342), .Z(n349) );
  GTECH_XOR2 U190 ( .A(cin), .B(n353), .Z(sum[0]) );
  GTECH_OAI21 U191 ( .A(n354), .B(n355), .C(n336), .Z(cout) );
  GTECH_OR3 U192 ( .A(n333), .B(n329), .C(n315), .Z(n336) );
  GTECH_AND2 U193 ( .A(b[12]), .B(a[12]), .Z(n329) );
  GTECH_NOT U194 ( .A(n315), .Z(n355) );
  GTECH_MUX2 U195 ( .A(n356), .B(n271), .S(n265), .Z(n315) );
  GTECH_NOT U196 ( .A(n268), .Z(n265) );
  GTECH_MUX2 U197 ( .A(n293), .B(n357), .S(n274), .Z(n268) );
  GTECH_MUX2 U198 ( .A(n353), .B(n358), .S(cin), .Z(n274) );
  GTECH_OA21 U199 ( .A(a[3]), .B(n297), .C(n359), .Z(n358) );
  GTECH_AO21 U200 ( .A(n297), .B(a[3]), .C(b[3]), .Z(n359) );
  GTECH_AO21 U201 ( .A(n299), .B(n305), .C(n301), .Z(n297) );
  GTECH_AND2 U202 ( .A(a[2]), .B(b[2]), .Z(n301) );
  GTECH_AO21 U203 ( .A(n312), .B(n306), .C(n308), .Z(n305) );
  GTECH_AND2 U204 ( .A(b[1]), .B(a[1]), .Z(n308) );
  GTECH_OR2 U205 ( .A(b[1]), .B(a[1]), .Z(n306) );
  GTECH_OR2 U206 ( .A(b[2]), .B(a[2]), .Z(n299) );
  GTECH_AND_NOT U207 ( .A(n312), .B(n307), .Z(n353) );
  GTECH_AND2 U208 ( .A(b[0]), .B(a[0]), .Z(n307) );
  GTECH_OR2 U209 ( .A(a[0]), .B(b[0]), .Z(n312) );
  GTECH_OAI21 U210 ( .A(n360), .B(n361), .C(n362), .Z(n357) );
  GTECH_OAI21 U211 ( .A(a[7]), .B(n276), .C(b[7]), .Z(n362) );
  GTECH_NOT U212 ( .A(n360), .Z(n276) );
  GTECH_NOT U213 ( .A(a[7]), .Z(n361) );
  GTECH_OA21 U214 ( .A(n285), .B(n278), .C(n280), .Z(n360) );
  GTECH_NAND2 U215 ( .A(b[6]), .B(a[6]), .Z(n280) );
  GTECH_NOR2 U216 ( .A(a[6]), .B(b[6]), .Z(n278) );
  GTECH_NOT U217 ( .A(n363), .Z(n285) );
  GTECH_AO21 U218 ( .A(n292), .B(n286), .C(n288), .Z(n363) );
  GTECH_AND2 U219 ( .A(b[5]), .B(a[5]), .Z(n288) );
  GTECH_OR2 U220 ( .A(b[5]), .B(a[5]), .Z(n286) );
  GTECH_AND_NOT U221 ( .A(n292), .B(n287), .Z(n293) );
  GTECH_AND2 U222 ( .A(b[4]), .B(a[4]), .Z(n287) );
  GTECH_OR2 U223 ( .A(a[4]), .B(b[4]), .Z(n292) );
  GTECH_XNOR2 U224 ( .A(n266), .B(b[8]), .Z(n271) );
  GTECH_NOT U225 ( .A(a[8]), .Z(n266) );
  GTECH_OA21 U226 ( .A(a[11]), .B(n346), .C(n364), .Z(n356) );
  GTECH_AO21 U227 ( .A(n346), .B(a[11]), .C(b[11]), .Z(n364) );
  GTECH_NAND2 U228 ( .A(n365), .B(n342), .Z(n346) );
  GTECH_NAND2 U229 ( .A(a[10]), .B(b[10]), .Z(n342) );
  GTECH_AO21 U230 ( .A(n344), .B(n343), .C(n352), .Z(n365) );
  GTECH_AND_NOT U231 ( .A(n366), .B(n351), .Z(n352) );
  GTECH_AND2 U232 ( .A(b[9]), .B(a[9]), .Z(n351) );
  GTECH_OAI21 U233 ( .A(b[8]), .B(a[8]), .C(n270), .Z(n366) );
  GTECH_OR2 U234 ( .A(b[9]), .B(a[9]), .Z(n270) );
  GTECH_NOT U235 ( .A(b[10]), .Z(n343) );
  GTECH_NOT U236 ( .A(a[10]), .Z(n344) );
  GTECH_OA21 U237 ( .A(n317), .B(n367), .C(n368), .Z(n354) );
  GTECH_OAI21 U238 ( .A(a[15]), .B(n369), .C(b[15]), .Z(n368) );
  GTECH_NOT U239 ( .A(a[15]), .Z(n367) );
  GTECH_NOT U240 ( .A(n369), .Z(n317) );
  GTECH_NAND2 U241 ( .A(n370), .B(n320), .Z(n369) );
  GTECH_NAND2 U242 ( .A(a[14]), .B(b[14]), .Z(n320) );
  GTECH_AO21 U243 ( .A(n322), .B(n321), .C(n327), .Z(n370) );
  GTECH_AOI2N2 U244 ( .A(a[13]), .B(b[13]), .C(n330), .D(n333), .Z(n327) );
  GTECH_NOR2 U245 ( .A(a[12]), .B(b[12]), .Z(n333) );
  GTECH_NOR2 U246 ( .A(a[13]), .B(b[13]), .Z(n330) );
  GTECH_NOT U247 ( .A(b[14]), .Z(n321) );
  GTECH_NOT U248 ( .A(a[14]), .Z(n322) );
endmodule

