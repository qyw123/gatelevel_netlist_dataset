
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_XOR2 U75 ( .A(n83), .B(n84), .Z(N155) );
  GTECH_AND2 U76 ( .A(n85), .B(n86), .Z(n84) );
  GTECH_OAI22 U77 ( .A(n87), .B(n88), .C(n89), .D(n90), .Z(n83) );
  GTECH_NOT U78 ( .A(n91), .Z(n90) );
  GTECH_XOR2 U79 ( .A(n85), .B(n86), .Z(N154) );
  GTECH_NOT U80 ( .A(n92), .Z(n86) );
  GTECH_XOR2 U81 ( .A(n91), .B(n89), .Z(n92) );
  GTECH_OA21 U82 ( .A(n93), .B(n94), .C(n95), .Z(n89) );
  GTECH_AO21 U83 ( .A(n94), .B(n93), .C(n96), .Z(n95) );
  GTECH_NOT U84 ( .A(n97), .Z(n94) );
  GTECH_XOR2 U85 ( .A(n88), .B(n87), .Z(n91) );
  GTECH_AOI2N2 U86 ( .A(n98), .B(n99), .C(n100), .D(n101), .Z(n87) );
  GTECH_NAND2 U87 ( .A(n100), .B(n101), .Z(n99) );
  GTECH_NAND2 U88 ( .A(I_b[7]), .B(I_a[7]), .Z(n88) );
  GTECH_NOT U89 ( .A(n102), .Z(n85) );
  GTECH_NAND2 U90 ( .A(n103), .B(n104), .Z(n102) );
  GTECH_XOR2 U91 ( .A(n104), .B(n103), .Z(N153) );
  GTECH_NOT U92 ( .A(n105), .Z(n103) );
  GTECH_XOR3 U93 ( .A(n106), .B(n96), .C(n97), .Z(n105) );
  GTECH_XOR3 U94 ( .A(n107), .B(n108), .C(n98), .Z(n97) );
  GTECH_OAI2N2 U95 ( .A(n109), .B(n110), .C(n111), .D(n112), .Z(n98) );
  GTECH_NAND2 U96 ( .A(n109), .B(n110), .Z(n112) );
  GTECH_NOT U97 ( .A(n101), .Z(n108) );
  GTECH_NAND2 U98 ( .A(I_a[7]), .B(I_b[6]), .Z(n101) );
  GTECH_NOT U99 ( .A(n100), .Z(n107) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n100) );
  GTECH_OA21 U101 ( .A(n113), .B(n114), .C(n115), .Z(n96) );
  GTECH_AO21 U102 ( .A(n113), .B(n114), .C(n116), .Z(n115) );
  GTECH_NOT U103 ( .A(n117), .Z(n113) );
  GTECH_NOT U104 ( .A(n93), .Z(n106) );
  GTECH_NAND2 U105 ( .A(I_a[7]), .B(n118), .Z(n93) );
  GTECH_NOT U106 ( .A(n119), .Z(n104) );
  GTECH_NAND2 U107 ( .A(n120), .B(n121), .Z(n119) );
  GTECH_XOR2 U108 ( .A(n122), .B(n123), .Z(N152) );
  GTECH_NOT U109 ( .A(n120), .Z(n123) );
  GTECH_XOR3 U110 ( .A(n116), .B(n114), .C(n117), .Z(n120) );
  GTECH_XOR2 U111 ( .A(n124), .B(n118), .Z(n117) );
  GTECH_OAI2N2 U112 ( .A(n125), .B(n126), .C(n127), .D(n128), .Z(n118) );
  GTECH_NAND2 U113 ( .A(n125), .B(n126), .Z(n128) );
  GTECH_AND2 U114 ( .A(I_a[7]), .B(I_b[5]), .Z(n124) );
  GTECH_NOT U115 ( .A(n129), .Z(n114) );
  GTECH_XOR3 U116 ( .A(n130), .B(n131), .C(n111), .Z(n129) );
  GTECH_OAI2N2 U117 ( .A(n132), .B(n133), .C(n134), .D(n135), .Z(n111) );
  GTECH_NAND2 U118 ( .A(n132), .B(n133), .Z(n135) );
  GTECH_NOT U119 ( .A(n110), .Z(n131) );
  GTECH_NAND2 U120 ( .A(I_b[6]), .B(I_a[6]), .Z(n110) );
  GTECH_NOT U121 ( .A(n109), .Z(n130) );
  GTECH_NAND2 U122 ( .A(I_b[7]), .B(I_a[5]), .Z(n109) );
  GTECH_OA21 U123 ( .A(n136), .B(n137), .C(n138), .Z(n116) );
  GTECH_AO21 U124 ( .A(n136), .B(n137), .C(n139), .Z(n138) );
  GTECH_NOT U125 ( .A(n140), .Z(n136) );
  GTECH_NOT U126 ( .A(n121), .Z(n122) );
  GTECH_OAI22 U127 ( .A(n141), .B(n142), .C(n143), .D(n144), .Z(n121) );
  GTECH_AND2 U128 ( .A(n141), .B(n142), .Z(n144) );
  GTECH_NOT U129 ( .A(n145), .Z(n142) );
  GTECH_XOR3 U130 ( .A(n143), .B(n141), .C(n145), .Z(N151) );
  GTECH_XOR3 U131 ( .A(n139), .B(n137), .C(n140), .Z(n145) );
  GTECH_XOR3 U132 ( .A(n146), .B(n147), .C(n127), .Z(n140) );
  GTECH_OAI2N2 U133 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n127) );
  GTECH_NAND2 U134 ( .A(n148), .B(n149), .Z(n151) );
  GTECH_NOT U135 ( .A(n126), .Z(n147) );
  GTECH_NAND2 U136 ( .A(I_a[7]), .B(I_b[4]), .Z(n126) );
  GTECH_NOT U137 ( .A(n125), .Z(n146) );
  GTECH_NAND2 U138 ( .A(I_a[6]), .B(I_b[5]), .Z(n125) );
  GTECH_NOT U139 ( .A(n152), .Z(n137) );
  GTECH_XOR3 U140 ( .A(n153), .B(n154), .C(n134), .Z(n152) );
  GTECH_OAI2N2 U141 ( .A(n155), .B(n156), .C(n157), .D(n158), .Z(n134) );
  GTECH_NAND2 U142 ( .A(n155), .B(n156), .Z(n158) );
  GTECH_NOT U143 ( .A(n133), .Z(n154) );
  GTECH_NAND2 U144 ( .A(I_b[6]), .B(I_a[5]), .Z(n133) );
  GTECH_NOT U145 ( .A(n132), .Z(n153) );
  GTECH_NAND2 U146 ( .A(I_b[7]), .B(I_a[4]), .Z(n132) );
  GTECH_OA21 U147 ( .A(n159), .B(n160), .C(n161), .Z(n139) );
  GTECH_AO21 U148 ( .A(n159), .B(n160), .C(n162), .Z(n161) );
  GTECH_NOT U149 ( .A(n163), .Z(n159) );
  GTECH_NOT U150 ( .A(n164), .Z(n141) );
  GTECH_OAI22 U151 ( .A(n165), .B(n166), .C(n167), .D(n168), .Z(n164) );
  GTECH_NOT U152 ( .A(I_a[7]), .Z(n167) );
  GTECH_OA21 U153 ( .A(n169), .B(n170), .C(n171), .Z(n143) );
  GTECH_AO21 U154 ( .A(n169), .B(n170), .C(n172), .Z(n171) );
  GTECH_NOT U155 ( .A(n173), .Z(n169) );
  GTECH_XOR3 U156 ( .A(n172), .B(n170), .C(n173), .Z(N150) );
  GTECH_XOR3 U157 ( .A(n162), .B(n160), .C(n163), .Z(n173) );
  GTECH_XOR3 U158 ( .A(n174), .B(n175), .C(n150), .Z(n163) );
  GTECH_OAI2N2 U159 ( .A(n176), .B(n177), .C(n178), .D(n179), .Z(n150) );
  GTECH_NAND2 U160 ( .A(n176), .B(n177), .Z(n179) );
  GTECH_NOT U161 ( .A(n149), .Z(n175) );
  GTECH_NAND2 U162 ( .A(I_a[6]), .B(I_b[4]), .Z(n149) );
  GTECH_NOT U163 ( .A(n148), .Z(n174) );
  GTECH_NAND2 U164 ( .A(I_b[5]), .B(I_a[5]), .Z(n148) );
  GTECH_NOT U165 ( .A(n180), .Z(n160) );
  GTECH_XOR3 U166 ( .A(n181), .B(n182), .C(n157), .Z(n180) );
  GTECH_OAI2N2 U167 ( .A(n183), .B(n184), .C(n185), .D(n186), .Z(n157) );
  GTECH_NAND2 U168 ( .A(n183), .B(n184), .Z(n186) );
  GTECH_NOT U169 ( .A(n156), .Z(n182) );
  GTECH_NAND2 U170 ( .A(I_b[6]), .B(I_a[4]), .Z(n156) );
  GTECH_NOT U171 ( .A(n155), .Z(n181) );
  GTECH_NAND2 U172 ( .A(I_b[7]), .B(I_a[3]), .Z(n155) );
  GTECH_OA21 U173 ( .A(n187), .B(n188), .C(n189), .Z(n162) );
  GTECH_AO21 U174 ( .A(n187), .B(n188), .C(n190), .Z(n189) );
  GTECH_NOT U175 ( .A(n191), .Z(n187) );
  GTECH_NOT U176 ( .A(n192), .Z(n170) );
  GTECH_XOR2 U177 ( .A(n166), .B(n165), .Z(n192) );
  GTECH_OA21 U178 ( .A(n193), .B(n194), .C(n195), .Z(n165) );
  GTECH_AO21 U179 ( .A(n193), .B(n194), .C(n196), .Z(n195) );
  GTECH_XOR2 U180 ( .A(n197), .B(n168), .Z(n166) );
  GTECH_OAI2N2 U181 ( .A(n198), .B(n199), .C(n200), .D(n201), .Z(n168) );
  GTECH_NAND2 U182 ( .A(n199), .B(n198), .Z(n201) );
  GTECH_AND2 U183 ( .A(I_a[7]), .B(I_b[3]), .Z(n197) );
  GTECH_OA21 U184 ( .A(n202), .B(n203), .C(n204), .Z(n172) );
  GTECH_AO21 U185 ( .A(n202), .B(n203), .C(n205), .Z(n204) );
  GTECH_NOT U186 ( .A(n206), .Z(n202) );
  GTECH_XOR3 U187 ( .A(n205), .B(n203), .C(n206), .Z(N149) );
  GTECH_XOR3 U188 ( .A(n190), .B(n188), .C(n191), .Z(n206) );
  GTECH_XOR3 U189 ( .A(n207), .B(n208), .C(n178), .Z(n191) );
  GTECH_OAI2N2 U190 ( .A(n209), .B(n210), .C(n211), .D(n212), .Z(n178) );
  GTECH_NAND2 U191 ( .A(n209), .B(n210), .Z(n212) );
  GTECH_NOT U192 ( .A(n177), .Z(n208) );
  GTECH_NAND2 U193 ( .A(I_a[5]), .B(I_b[4]), .Z(n177) );
  GTECH_NOT U194 ( .A(n176), .Z(n207) );
  GTECH_NAND2 U195 ( .A(I_b[5]), .B(I_a[4]), .Z(n176) );
  GTECH_NOT U196 ( .A(n213), .Z(n188) );
  GTECH_XOR3 U197 ( .A(n214), .B(n215), .C(n185), .Z(n213) );
  GTECH_AO21 U198 ( .A(n216), .B(n217), .C(n218), .Z(n185) );
  GTECH_NOT U199 ( .A(n219), .Z(n218) );
  GTECH_NOT U200 ( .A(n184), .Z(n215) );
  GTECH_NAND2 U201 ( .A(I_b[6]), .B(I_a[3]), .Z(n184) );
  GTECH_NOT U202 ( .A(n183), .Z(n214) );
  GTECH_NAND2 U203 ( .A(I_b[7]), .B(I_a[2]), .Z(n183) );
  GTECH_OA21 U204 ( .A(n220), .B(n221), .C(n222), .Z(n190) );
  GTECH_AO21 U205 ( .A(n220), .B(n221), .C(n223), .Z(n222) );
  GTECH_NOT U206 ( .A(n224), .Z(n203) );
  GTECH_XOR3 U207 ( .A(n225), .B(n196), .C(n193), .Z(n224) );
  GTECH_XOR3 U208 ( .A(n198), .B(n199), .C(n200), .Z(n193) );
  GTECH_OAI22 U209 ( .A(n226), .B(n227), .C(n228), .D(n229), .Z(n200) );
  GTECH_AND2 U210 ( .A(n227), .B(n226), .Z(n228) );
  GTECH_NOT U211 ( .A(n230), .Z(n199) );
  GTECH_NAND2 U212 ( .A(I_a[7]), .B(I_b[2]), .Z(n230) );
  GTECH_NOT U213 ( .A(n231), .Z(n198) );
  GTECH_NAND2 U214 ( .A(I_a[6]), .B(I_b[3]), .Z(n231) );
  GTECH_OA21 U215 ( .A(n232), .B(n233), .C(n234), .Z(n196) );
  GTECH_AO21 U216 ( .A(n232), .B(n233), .C(n235), .Z(n234) );
  GTECH_NOT U217 ( .A(n236), .Z(n232) );
  GTECH_NOT U218 ( .A(n194), .Z(n225) );
  GTECH_NAND2 U219 ( .A(I_a[7]), .B(n237), .Z(n194) );
  GTECH_OA21 U220 ( .A(n238), .B(n239), .C(n240), .Z(n205) );
  GTECH_AO21 U221 ( .A(n238), .B(n239), .C(n241), .Z(n240) );
  GTECH_XOR3 U222 ( .A(n241), .B(n239), .C(n242), .Z(N148) );
  GTECH_NOT U223 ( .A(n238), .Z(n242) );
  GTECH_XOR3 U224 ( .A(n223), .B(n221), .C(n220), .Z(n238) );
  GTECH_XOR3 U225 ( .A(n217), .B(n216), .C(n219), .Z(n220) );
  GTECH_NAND3 U226 ( .A(I_b[7]), .B(I_a[0]), .C(n243), .Z(n219) );
  GTECH_NOT U227 ( .A(n244), .Z(n216) );
  GTECH_NAND2 U228 ( .A(I_b[6]), .B(I_a[2]), .Z(n244) );
  GTECH_NOT U229 ( .A(n245), .Z(n217) );
  GTECH_NAND2 U230 ( .A(I_b[7]), .B(I_a[1]), .Z(n245) );
  GTECH_NOT U231 ( .A(n246), .Z(n221) );
  GTECH_XOR3 U232 ( .A(n247), .B(n248), .C(n211), .Z(n246) );
  GTECH_OAI2N2 U233 ( .A(n249), .B(n250), .C(n251), .D(n252), .Z(n211) );
  GTECH_NAND2 U234 ( .A(n249), .B(n250), .Z(n252) );
  GTECH_NOT U235 ( .A(n210), .Z(n248) );
  GTECH_NAND2 U236 ( .A(I_b[4]), .B(I_a[4]), .Z(n210) );
  GTECH_NOT U237 ( .A(n209), .Z(n247) );
  GTECH_NAND2 U238 ( .A(I_b[5]), .B(I_a[3]), .Z(n209) );
  GTECH_OA21 U239 ( .A(n253), .B(n254), .C(n255), .Z(n223) );
  GTECH_AO21 U240 ( .A(n253), .B(n254), .C(n256), .Z(n255) );
  GTECH_NOT U241 ( .A(n257), .Z(n239) );
  GTECH_XOR3 U242 ( .A(n235), .B(n233), .C(n236), .Z(n257) );
  GTECH_XOR2 U243 ( .A(n258), .B(n237), .Z(n236) );
  GTECH_OAI2N2 U244 ( .A(n259), .B(n260), .C(n261), .D(n262), .Z(n237) );
  GTECH_NAND2 U245 ( .A(n259), .B(n260), .Z(n262) );
  GTECH_AND2 U246 ( .A(I_a[7]), .B(I_b[1]), .Z(n258) );
  GTECH_NOT U247 ( .A(n263), .Z(n233) );
  GTECH_XOR3 U248 ( .A(n226), .B(n227), .C(n229), .Z(n263) );
  GTECH_OAI2N2 U249 ( .A(n264), .B(n265), .C(n266), .D(n267), .Z(n229) );
  GTECH_NAND2 U250 ( .A(n264), .B(n265), .Z(n267) );
  GTECH_NOT U251 ( .A(n268), .Z(n227) );
  GTECH_NAND2 U252 ( .A(I_a[6]), .B(I_b[2]), .Z(n268) );
  GTECH_NOT U253 ( .A(n269), .Z(n226) );
  GTECH_NAND2 U254 ( .A(I_a[5]), .B(I_b[3]), .Z(n269) );
  GTECH_OA21 U255 ( .A(n270), .B(n271), .C(n272), .Z(n235) );
  GTECH_AO21 U256 ( .A(n270), .B(n271), .C(n273), .Z(n272) );
  GTECH_NOT U257 ( .A(n274), .Z(n270) );
  GTECH_OA21 U258 ( .A(n275), .B(n276), .C(n277), .Z(n241) );
  GTECH_AO21 U259 ( .A(n275), .B(n276), .C(n278), .Z(n277) );
  GTECH_NOT U260 ( .A(n279), .Z(n275) );
  GTECH_XOR3 U261 ( .A(n278), .B(n276), .C(n279), .Z(N147) );
  GTECH_XOR3 U262 ( .A(n280), .B(n254), .C(n253), .Z(n279) );
  GTECH_XOR2 U263 ( .A(n281), .B(n243), .Z(n253) );
  GTECH_NOT U264 ( .A(n282), .Z(n243) );
  GTECH_NAND2 U265 ( .A(I_b[6]), .B(I_a[1]), .Z(n282) );
  GTECH_NAND2 U266 ( .A(I_b[7]), .B(I_a[0]), .Z(n281) );
  GTECH_NOT U267 ( .A(n283), .Z(n254) );
  GTECH_XOR3 U268 ( .A(n284), .B(n285), .C(n251), .Z(n283) );
  GTECH_AO21 U269 ( .A(n286), .B(n287), .C(n288), .Z(n251) );
  GTECH_NOT U270 ( .A(n289), .Z(n288) );
  GTECH_NOT U271 ( .A(n250), .Z(n285) );
  GTECH_NAND2 U272 ( .A(I_b[4]), .B(I_a[3]), .Z(n250) );
  GTECH_NOT U273 ( .A(n249), .Z(n284) );
  GTECH_NAND2 U274 ( .A(I_b[5]), .B(I_a[2]), .Z(n249) );
  GTECH_NOT U275 ( .A(n256), .Z(n280) );
  GTECH_NAND3 U276 ( .A(I_a[0]), .B(n290), .C(I_b[6]), .Z(n256) );
  GTECH_NOT U277 ( .A(n291), .Z(n290) );
  GTECH_NOT U278 ( .A(n292), .Z(n276) );
  GTECH_XOR3 U279 ( .A(n273), .B(n271), .C(n274), .Z(n292) );
  GTECH_XOR3 U280 ( .A(n293), .B(n294), .C(n261), .Z(n274) );
  GTECH_OAI2N2 U281 ( .A(n295), .B(n296), .C(n297), .D(n298), .Z(n261) );
  GTECH_NAND2 U282 ( .A(n295), .B(n296), .Z(n298) );
  GTECH_NOT U283 ( .A(n260), .Z(n294) );
  GTECH_NAND2 U284 ( .A(I_a[7]), .B(I_b[0]), .Z(n260) );
  GTECH_NOT U285 ( .A(n259), .Z(n293) );
  GTECH_NAND2 U286 ( .A(I_a[6]), .B(I_b[1]), .Z(n259) );
  GTECH_NOT U287 ( .A(n299), .Z(n271) );
  GTECH_XOR3 U288 ( .A(n300), .B(n301), .C(n266), .Z(n299) );
  GTECH_OAI2N2 U289 ( .A(n302), .B(n303), .C(n304), .D(n305), .Z(n266) );
  GTECH_NAND2 U290 ( .A(n302), .B(n303), .Z(n305) );
  GTECH_NOT U291 ( .A(n265), .Z(n301) );
  GTECH_NAND2 U292 ( .A(I_a[5]), .B(I_b[2]), .Z(n265) );
  GTECH_NOT U293 ( .A(n264), .Z(n300) );
  GTECH_NAND2 U294 ( .A(I_a[4]), .B(I_b[3]), .Z(n264) );
  GTECH_OA21 U295 ( .A(n306), .B(n307), .C(n308), .Z(n273) );
  GTECH_AO21 U296 ( .A(n306), .B(n307), .C(n309), .Z(n308) );
  GTECH_NOT U297 ( .A(n310), .Z(n306) );
  GTECH_OA21 U298 ( .A(n311), .B(n312), .C(n313), .Z(n278) );
  GTECH_AO21 U299 ( .A(n311), .B(n312), .C(n314), .Z(n313) );
  GTECH_XOR3 U300 ( .A(n314), .B(n312), .C(n315), .Z(N146) );
  GTECH_NOT U301 ( .A(n311), .Z(n315) );
  GTECH_XOR2 U302 ( .A(n291), .B(n316), .Z(n311) );
  GTECH_AND2 U303 ( .A(I_b[6]), .B(I_a[0]), .Z(n316) );
  GTECH_XOR3 U304 ( .A(n287), .B(n286), .C(n289), .Z(n291) );
  GTECH_NAND3 U305 ( .A(I_b[5]), .B(I_a[0]), .C(n317), .Z(n289) );
  GTECH_NOT U306 ( .A(n318), .Z(n286) );
  GTECH_NAND2 U307 ( .A(I_b[4]), .B(I_a[2]), .Z(n318) );
  GTECH_NOT U308 ( .A(n319), .Z(n287) );
  GTECH_NAND2 U309 ( .A(I_b[5]), .B(I_a[1]), .Z(n319) );
  GTECH_NOT U310 ( .A(n320), .Z(n312) );
  GTECH_XOR3 U311 ( .A(n309), .B(n307), .C(n310), .Z(n320) );
  GTECH_XOR3 U312 ( .A(n321), .B(n322), .C(n297), .Z(n310) );
  GTECH_OAI2N2 U313 ( .A(n323), .B(n324), .C(n325), .D(n326), .Z(n297) );
  GTECH_NAND2 U314 ( .A(n323), .B(n324), .Z(n326) );
  GTECH_NOT U315 ( .A(n296), .Z(n322) );
  GTECH_NAND2 U316 ( .A(I_a[6]), .B(I_b[0]), .Z(n296) );
  GTECH_NOT U317 ( .A(n295), .Z(n321) );
  GTECH_NAND2 U318 ( .A(I_a[5]), .B(I_b[1]), .Z(n295) );
  GTECH_NOT U319 ( .A(n327), .Z(n307) );
  GTECH_XOR3 U320 ( .A(n328), .B(n329), .C(n304), .Z(n327) );
  GTECH_OAI2N2 U321 ( .A(n330), .B(n331), .C(n332), .D(n333), .Z(n304) );
  GTECH_NAND2 U322 ( .A(n330), .B(n331), .Z(n333) );
  GTECH_NOT U323 ( .A(n303), .Z(n329) );
  GTECH_NAND2 U324 ( .A(I_a[4]), .B(I_b[2]), .Z(n303) );
  GTECH_NOT U325 ( .A(n302), .Z(n328) );
  GTECH_NAND2 U326 ( .A(I_a[3]), .B(I_b[3]), .Z(n302) );
  GTECH_OA21 U327 ( .A(n334), .B(n335), .C(n336), .Z(n309) );
  GTECH_AO21 U328 ( .A(n334), .B(n335), .C(n337), .Z(n336) );
  GTECH_NOT U329 ( .A(n338), .Z(n334) );
  GTECH_OA21 U330 ( .A(n339), .B(n340), .C(n341), .Z(n314) );
  GTECH_AO21 U331 ( .A(n339), .B(n340), .C(n342), .Z(n341) );
  GTECH_XOR3 U332 ( .A(n343), .B(n340), .C(n339), .Z(N145) );
  GTECH_XOR2 U333 ( .A(n344), .B(n317), .Z(n339) );
  GTECH_NOT U334 ( .A(n345), .Z(n317) );
  GTECH_NAND2 U335 ( .A(I_b[4]), .B(I_a[1]), .Z(n345) );
  GTECH_NAND2 U336 ( .A(I_b[5]), .B(I_a[0]), .Z(n344) );
  GTECH_NOT U337 ( .A(n346), .Z(n340) );
  GTECH_XOR3 U338 ( .A(n337), .B(n335), .C(n338), .Z(n346) );
  GTECH_XOR3 U339 ( .A(n347), .B(n348), .C(n325), .Z(n338) );
  GTECH_OAI2N2 U340 ( .A(n349), .B(n350), .C(n351), .D(n352), .Z(n325) );
  GTECH_NAND2 U341 ( .A(n349), .B(n350), .Z(n352) );
  GTECH_NOT U342 ( .A(n324), .Z(n348) );
  GTECH_NAND2 U343 ( .A(I_a[5]), .B(I_b[0]), .Z(n324) );
  GTECH_NOT U344 ( .A(n323), .Z(n347) );
  GTECH_NAND2 U345 ( .A(I_a[4]), .B(I_b[1]), .Z(n323) );
  GTECH_NOT U346 ( .A(n353), .Z(n335) );
  GTECH_XOR3 U347 ( .A(n354), .B(n355), .C(n332), .Z(n353) );
  GTECH_AO21 U348 ( .A(n356), .B(n357), .C(n358), .Z(n332) );
  GTECH_NOT U349 ( .A(n359), .Z(n358) );
  GTECH_NOT U350 ( .A(n331), .Z(n355) );
  GTECH_NAND2 U351 ( .A(I_a[3]), .B(I_b[2]), .Z(n331) );
  GTECH_NOT U352 ( .A(n330), .Z(n354) );
  GTECH_NAND2 U353 ( .A(I_a[2]), .B(I_b[3]), .Z(n330) );
  GTECH_OA21 U354 ( .A(n360), .B(n361), .C(n362), .Z(n337) );
  GTECH_AO21 U355 ( .A(n360), .B(n361), .C(n363), .Z(n362) );
  GTECH_NOT U356 ( .A(n342), .Z(n343) );
  GTECH_NAND3 U357 ( .A(I_a[0]), .B(n364), .C(I_b[4]), .Z(n342) );
  GTECH_XOR2 U358 ( .A(n365), .B(n364), .Z(N144) );
  GTECH_NOT U359 ( .A(n366), .Z(n364) );
  GTECH_XOR3 U360 ( .A(n363), .B(n361), .C(n360), .Z(n366) );
  GTECH_XOR3 U361 ( .A(n357), .B(n356), .C(n359), .Z(n360) );
  GTECH_NAND3 U362 ( .A(I_a[0]), .B(n367), .C(I_b[3]), .Z(n359) );
  GTECH_NOT U363 ( .A(n368), .Z(n356) );
  GTECH_NAND2 U364 ( .A(I_a[2]), .B(I_b[2]), .Z(n368) );
  GTECH_NOT U365 ( .A(n369), .Z(n357) );
  GTECH_NAND2 U366 ( .A(I_b[3]), .B(I_a[1]), .Z(n369) );
  GTECH_NOT U367 ( .A(n370), .Z(n361) );
  GTECH_XOR3 U368 ( .A(n371), .B(n372), .C(n351), .Z(n370) );
  GTECH_OAI2N2 U369 ( .A(n373), .B(n374), .C(n375), .D(n376), .Z(n351) );
  GTECH_NAND2 U370 ( .A(n373), .B(n374), .Z(n376) );
  GTECH_NOT U371 ( .A(n350), .Z(n372) );
  GTECH_NAND2 U372 ( .A(I_a[4]), .B(I_b[0]), .Z(n350) );
  GTECH_NOT U373 ( .A(n349), .Z(n371) );
  GTECH_NAND2 U374 ( .A(I_a[3]), .B(I_b[1]), .Z(n349) );
  GTECH_OA21 U375 ( .A(n377), .B(n378), .C(n379), .Z(n363) );
  GTECH_AO21 U376 ( .A(n377), .B(n378), .C(n380), .Z(n379) );
  GTECH_AND2 U377 ( .A(I_b[4]), .B(I_a[0]), .Z(n365) );
  GTECH_XOR3 U378 ( .A(n381), .B(n378), .C(n377), .Z(N143) );
  GTECH_XOR2 U379 ( .A(n382), .B(n367), .Z(n377) );
  GTECH_NOT U380 ( .A(n383), .Z(n367) );
  GTECH_NAND2 U381 ( .A(I_b[2]), .B(I_a[1]), .Z(n383) );
  GTECH_NAND2 U382 ( .A(I_b[3]), .B(I_a[0]), .Z(n382) );
  GTECH_NOT U383 ( .A(n384), .Z(n378) );
  GTECH_XOR3 U384 ( .A(n385), .B(n386), .C(n375), .Z(n384) );
  GTECH_AO21 U385 ( .A(n387), .B(n388), .C(n389), .Z(n375) );
  GTECH_NOT U386 ( .A(n390), .Z(n389) );
  GTECH_NOT U387 ( .A(n374), .Z(n386) );
  GTECH_NAND2 U388 ( .A(I_a[3]), .B(I_b[0]), .Z(n374) );
  GTECH_NOT U389 ( .A(n373), .Z(n385) );
  GTECH_NAND2 U390 ( .A(I_b[1]), .B(I_a[2]), .Z(n373) );
  GTECH_NOT U391 ( .A(n380), .Z(n381) );
  GTECH_NAND3 U392 ( .A(I_b[2]), .B(n391), .C(I_a[0]), .Z(n380) );
  GTECH_XOR2 U393 ( .A(n392), .B(n391), .Z(N142) );
  GTECH_NOT U394 ( .A(n393), .Z(n391) );
  GTECH_XOR3 U395 ( .A(n388), .B(n387), .C(n390), .Z(n393) );
  GTECH_NAND3 U396 ( .A(n394), .B(I_a[0]), .C(I_b[1]), .Z(n390) );
  GTECH_NOT U397 ( .A(n395), .Z(n387) );
  GTECH_NAND2 U398 ( .A(I_b[0]), .B(I_a[2]), .Z(n395) );
  GTECH_NOT U399 ( .A(n396), .Z(n388) );
  GTECH_NAND2 U400 ( .A(I_b[1]), .B(I_a[1]), .Z(n396) );
  GTECH_AND2 U401 ( .A(I_a[0]), .B(I_b[2]), .Z(n392) );
  GTECH_XOR2 U402 ( .A(n394), .B(n397), .Z(N141) );
  GTECH_AND2 U403 ( .A(I_b[1]), .B(I_a[0]), .Z(n397) );
  GTECH_NOT U404 ( .A(n398), .Z(n394) );
  GTECH_NAND2 U405 ( .A(I_b[0]), .B(I_a[1]), .Z(n398) );
  GTECH_AND2 U406 ( .A(I_b[0]), .B(I_a[0]), .Z(N140) );
endmodule

