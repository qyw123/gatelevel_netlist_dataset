
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373;

  GTECH_MUX2 U127 ( .A(n266), .B(n267), .S(n268), .Z(sum[9]) );
  GTECH_XNOR2 U128 ( .A(n269), .B(n270), .Z(n267) );
  GTECH_XOR2 U129 ( .A(n270), .B(n271), .Z(n266) );
  GTECH_OAI21 U130 ( .A(b[9]), .B(a[9]), .C(n272), .Z(n270) );
  GTECH_XNOR2 U131 ( .A(n273), .B(n274), .Z(sum[8]) );
  GTECH_MUX2 U132 ( .A(n275), .B(n276), .S(n277), .Z(sum[7]) );
  GTECH_XOR2 U133 ( .A(n278), .B(n279), .Z(n276) );
  GTECH_OA21 U134 ( .A(n280), .B(n281), .C(n282), .Z(n279) );
  GTECH_XNOR2 U135 ( .A(n278), .B(n283), .Z(n275) );
  GTECH_XNOR2 U136 ( .A(a[7]), .B(b[7]), .Z(n278) );
  GTECH_MUX2 U137 ( .A(n284), .B(n285), .S(n286), .Z(sum[6]) );
  GTECH_XNOR2 U138 ( .A(n287), .B(n288), .Z(n285) );
  GTECH_XNOR2 U139 ( .A(n281), .B(n287), .Z(n284) );
  GTECH_NOR2 U140 ( .A(n280), .B(n289), .Z(n287) );
  GTECH_AOI21 U141 ( .A(b[4]), .B(n290), .C(n291), .Z(n281) );
  GTECH_AND2 U142 ( .A(n292), .B(a[4]), .Z(n290) );
  GTECH_XNOR2 U143 ( .A(n293), .B(n294), .Z(sum[5]) );
  GTECH_OR_NOT U144 ( .A(n291), .B(n292), .Z(n294) );
  GTECH_AND2 U145 ( .A(n295), .B(n296), .Z(n293) );
  GTECH_AO21 U146 ( .A(a[4]), .B(b[4]), .C(n286), .Z(n296) );
  GTECH_XNOR2 U147 ( .A(n277), .B(n297), .Z(sum[4]) );
  GTECH_MUX2 U148 ( .A(n298), .B(n299), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U149 ( .A(n300), .B(n301), .Z(n299) );
  GTECH_XOR2 U150 ( .A(n300), .B(n302), .Z(n298) );
  GTECH_OA21 U151 ( .A(n303), .B(n304), .C(n305), .Z(n302) );
  GTECH_XNOR2 U152 ( .A(a[3]), .B(b[3]), .Z(n300) );
  GTECH_MUX2 U153 ( .A(n306), .B(n307), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U154 ( .A(n308), .B(n309), .Z(n307) );
  GTECH_XOR2 U155 ( .A(n304), .B(n308), .Z(n306) );
  GTECH_OR_NOT U156 ( .A(n303), .B(n305), .Z(n308) );
  GTECH_OA21 U157 ( .A(n310), .B(n311), .C(n312), .Z(n304) );
  GTECH_MUX2 U158 ( .A(n313), .B(n314), .S(n315), .Z(sum[1]) );
  GTECH_NOR2 U159 ( .A(n316), .B(n310), .Z(n315) );
  GTECH_AO21 U160 ( .A(n317), .B(n311), .C(n318), .Z(n314) );
  GTECH_OAI21 U161 ( .A(n318), .B(n317), .C(n311), .Z(n313) );
  GTECH_OR_NOT U162 ( .A(n319), .B(a[0]), .Z(n311) );
  GTECH_MUX2 U163 ( .A(n320), .B(n321), .S(n322), .Z(sum[15]) );
  GTECH_XOR2 U164 ( .A(n323), .B(n324), .Z(n321) );
  GTECH_AND2 U165 ( .A(n325), .B(n326), .Z(n324) );
  GTECH_OAI21 U166 ( .A(b[14]), .B(a[14]), .C(n327), .Z(n326) );
  GTECH_OA21 U167 ( .A(n328), .B(n329), .C(n330), .Z(n327) );
  GTECH_XNOR2 U168 ( .A(n323), .B(n331), .Z(n320) );
  GTECH_XNOR2 U169 ( .A(a[15]), .B(b[15]), .Z(n323) );
  GTECH_OAI21 U170 ( .A(n332), .B(n325), .C(n333), .Z(sum[14]) );
  GTECH_MUX2 U171 ( .A(n334), .B(n335), .S(b[14]), .Z(n333) );
  GTECH_OR_NOT U172 ( .A(a[14]), .B(n332), .Z(n335) );
  GTECH_XOR2 U173 ( .A(a[14]), .B(n332), .Z(n334) );
  GTECH_OA21 U174 ( .A(n336), .B(n322), .C(n337), .Z(n332) );
  GTECH_AOI21 U175 ( .A(n330), .B(n328), .C(n329), .Z(n337) );
  GTECH_MUX2 U176 ( .A(n338), .B(n339), .S(n322), .Z(sum[13]) );
  GTECH_XNOR2 U177 ( .A(n328), .B(n340), .Z(n339) );
  GTECH_XNOR2 U178 ( .A(n340), .B(n341), .Z(n338) );
  GTECH_OR_NOT U179 ( .A(n329), .B(n330), .Z(n340) );
  GTECH_OAI21 U180 ( .A(n342), .B(n322), .C(n343), .Z(sum[12]) );
  GTECH_AND2 U181 ( .A(n341), .B(n344), .Z(n342) );
  GTECH_MUX2 U182 ( .A(n345), .B(n346), .S(n268), .Z(sum[11]) );
  GTECH_XOR2 U183 ( .A(n347), .B(n348), .Z(n346) );
  GTECH_OA21 U184 ( .A(n349), .B(n350), .C(n351), .Z(n348) );
  GTECH_XNOR2 U185 ( .A(n347), .B(n352), .Z(n345) );
  GTECH_XNOR2 U186 ( .A(a[11]), .B(b[11]), .Z(n347) );
  GTECH_MUX2 U187 ( .A(n353), .B(n354), .S(n268), .Z(sum[10]) );
  GTECH_XNOR2 U188 ( .A(n350), .B(n355), .Z(n354) );
  GTECH_AOI21 U189 ( .A(n356), .B(n269), .C(n357), .Z(n350) );
  GTECH_NOT U190 ( .A(n358), .Z(n356) );
  GTECH_XNOR2 U191 ( .A(n355), .B(n359), .Z(n353) );
  GTECH_NOR2 U192 ( .A(n349), .B(n360), .Z(n355) );
  GTECH_XNOR2 U193 ( .A(n317), .B(n361), .Z(sum[0]) );
  GTECH_NOT U194 ( .A(cin), .Z(n317) );
  GTECH_OAI21 U195 ( .A(n362), .B(n322), .C(n343), .Z(cout) );
  GTECH_NAND3 U196 ( .A(n341), .B(n344), .C(n322), .Z(n343) );
  GTECH_NOT U197 ( .A(n328), .Z(n344) );
  GTECH_AND2 U198 ( .A(a[12]), .B(b[12]), .Z(n328) );
  GTECH_MUX2 U199 ( .A(n363), .B(n274), .S(n268), .Z(n322) );
  GTECH_NOT U200 ( .A(n273), .Z(n268) );
  GTECH_MUX2 U201 ( .A(n364), .B(n297), .S(n277), .Z(n273) );
  GTECH_NOT U202 ( .A(n286), .Z(n277) );
  GTECH_MUX2 U203 ( .A(n361), .B(n365), .S(cin), .Z(n286) );
  GTECH_OA21 U204 ( .A(a[3]), .B(n301), .C(n366), .Z(n365) );
  GTECH_AO21 U205 ( .A(n301), .B(a[3]), .C(b[3]), .Z(n366) );
  GTECH_OAI21 U206 ( .A(n309), .B(n303), .C(n305), .Z(n301) );
  GTECH_NOT U207 ( .A(n367), .Z(n305) );
  GTECH_AND2 U208 ( .A(a[2]), .B(b[2]), .Z(n367) );
  GTECH_NOR2 U209 ( .A(a[2]), .B(b[2]), .Z(n303) );
  GTECH_OA21 U210 ( .A(n310), .B(n318), .C(n312), .Z(n309) );
  GTECH_NOT U211 ( .A(n316), .Z(n312) );
  GTECH_AND2 U212 ( .A(a[1]), .B(b[1]), .Z(n316) );
  GTECH_NOR2 U213 ( .A(a[0]), .B(b[0]), .Z(n318) );
  GTECH_NOR2 U214 ( .A(a[1]), .B(b[1]), .Z(n310) );
  GTECH_XNOR2 U215 ( .A(a[0]), .B(n319), .Z(n361) );
  GTECH_NOT U216 ( .A(b[0]), .Z(n319) );
  GTECH_AOI21 U217 ( .A(a[4]), .B(b[4]), .C(n368), .Z(n297) );
  GTECH_OA21 U218 ( .A(a[7]), .B(n283), .C(n369), .Z(n364) );
  GTECH_AO21 U219 ( .A(n283), .B(a[7]), .C(b[7]), .Z(n369) );
  GTECH_OAI21 U220 ( .A(n288), .B(n280), .C(n282), .Z(n283) );
  GTECH_NOT U221 ( .A(n289), .Z(n282) );
  GTECH_AND2 U222 ( .A(a[6]), .B(b[6]), .Z(n289) );
  GTECH_NOR2 U223 ( .A(a[6]), .B(b[6]), .Z(n280) );
  GTECH_AOI21 U224 ( .A(n295), .B(n292), .C(n291), .Z(n288) );
  GTECH_AND2 U225 ( .A(a[5]), .B(b[5]), .Z(n291) );
  GTECH_OR2 U226 ( .A(a[5]), .B(b[5]), .Z(n292) );
  GTECH_NOT U227 ( .A(n368), .Z(n295) );
  GTECH_NOR2 U228 ( .A(b[4]), .B(a[4]), .Z(n368) );
  GTECH_OR2 U229 ( .A(n271), .B(n269), .Z(n274) );
  GTECH_AND2 U230 ( .A(a[8]), .B(b[8]), .Z(n269) );
  GTECH_AOI21 U231 ( .A(n352), .B(a[11]), .C(n370), .Z(n363) );
  GTECH_OA21 U232 ( .A(a[11]), .B(n352), .C(b[11]), .Z(n370) );
  GTECH_OAI21 U233 ( .A(n359), .B(n349), .C(n351), .Z(n352) );
  GTECH_NOT U234 ( .A(n360), .Z(n351) );
  GTECH_AND2 U235 ( .A(a[10]), .B(b[10]), .Z(n360) );
  GTECH_NOR2 U236 ( .A(a[10]), .B(b[10]), .Z(n349) );
  GTECH_OA21 U237 ( .A(n358), .B(n271), .C(n272), .Z(n359) );
  GTECH_NOT U238 ( .A(n357), .Z(n272) );
  GTECH_AND2 U239 ( .A(a[9]), .B(b[9]), .Z(n357) );
  GTECH_NOR2 U240 ( .A(a[8]), .B(b[8]), .Z(n271) );
  GTECH_NOR2 U241 ( .A(a[9]), .B(b[9]), .Z(n358) );
  GTECH_AOI21 U242 ( .A(n331), .B(a[15]), .C(n371), .Z(n362) );
  GTECH_OA21 U243 ( .A(a[15]), .B(n331), .C(b[15]), .Z(n371) );
  GTECH_OAI21 U244 ( .A(n336), .B(n372), .C(n325), .Z(n331) );
  GTECH_NOT U245 ( .A(n373), .Z(n325) );
  GTECH_AND2 U246 ( .A(a[14]), .B(b[14]), .Z(n373) );
  GTECH_NOR2 U247 ( .A(a[14]), .B(b[14]), .Z(n372) );
  GTECH_AOI21 U248 ( .A(n341), .B(n330), .C(n329), .Z(n336) );
  GTECH_AND2 U249 ( .A(a[13]), .B(b[13]), .Z(n329) );
  GTECH_OR2 U250 ( .A(a[13]), .B(b[13]), .Z(n330) );
  GTECH_OR2 U251 ( .A(b[12]), .B(a[12]), .Z(n341) );
endmodule

