
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_OAI21 U75 ( .A(n83), .B(n84), .C(n85), .Z(N155) );
  GTECH_OA22 U76 ( .A(n86), .B(n87), .C(n88), .D(n89), .Z(n85) );
  GTECH_XNOR2 U77 ( .A(n90), .B(n83), .Z(N154) );
  GTECH_XNOR2 U78 ( .A(n86), .B(n87), .Z(n83) );
  GTECH_NOT U79 ( .A(n91), .Z(n87) );
  GTECH_XNOR2 U80 ( .A(n88), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n89), .Z(n92) );
  GTECH_NAND2 U82 ( .A(I_b[7]), .B(I_a[7]), .Z(n89) );
  GTECH_AND2 U83 ( .A(n93), .B(n94), .Z(n88) );
  GTECH_OR_NOT U84 ( .A(n95), .B(n96), .Z(n94) );
  GTECH_OAI21 U85 ( .A(n97), .B(n96), .C(n98), .Z(n93) );
  GTECH_AOI2N2 U86 ( .A(n99), .B(n100), .C(n101), .D(n102), .Z(n86) );
  GTECH_NAND2 U87 ( .A(n101), .B(n102), .Z(n100) );
  GTECH_NOT U88 ( .A(n84), .Z(n90) );
  GTECH_NAND2 U89 ( .A(n103), .B(n104), .Z(n84) );
  GTECH_NOT U90 ( .A(n105), .Z(n103) );
  GTECH_XNOR2 U91 ( .A(n104), .B(n105), .Z(N153) );
  GTECH_XOR3 U92 ( .A(n106), .B(n101), .C(n99), .Z(n105) );
  GTECH_XOR3 U93 ( .A(n97), .B(n98), .C(n96), .Z(n99) );
  GTECH_OAI21 U94 ( .A(n107), .B(n108), .C(n109), .Z(n96) );
  GTECH_OAI21 U95 ( .A(n110), .B(n111), .C(n112), .Z(n109) );
  GTECH_NOT U96 ( .A(n111), .Z(n107) );
  GTECH_NOT U97 ( .A(n113), .Z(n98) );
  GTECH_NAND2 U98 ( .A(I_b[7]), .B(I_a[6]), .Z(n113) );
  GTECH_NOT U99 ( .A(n95), .Z(n97) );
  GTECH_NAND2 U100 ( .A(I_a[7]), .B(I_b[6]), .Z(n95) );
  GTECH_ADD_ABC U101 ( .A(n114), .B(n115), .C(n116), .COUT(n101) );
  GTECH_NOT U102 ( .A(n117), .Z(n116) );
  GTECH_XNOR2 U103 ( .A(n118), .B(n119), .Z(n115) );
  GTECH_NAND2 U104 ( .A(I_a[7]), .B(I_b[5]), .Z(n119) );
  GTECH_NOT U105 ( .A(n102), .Z(n106) );
  GTECH_NAND2 U106 ( .A(I_a[7]), .B(n120), .Z(n102) );
  GTECH_NOT U107 ( .A(n121), .Z(n104) );
  GTECH_NAND2 U108 ( .A(n122), .B(n123), .Z(n121) );
  GTECH_NOT U109 ( .A(n124), .Z(n123) );
  GTECH_XNOR2 U110 ( .A(n124), .B(n122), .Z(N152) );
  GTECH_XOR4 U111 ( .A(n118), .B(n125), .C(n114), .D(n117), .Z(n122) );
  GTECH_XOR3 U112 ( .A(n110), .B(n112), .C(n111), .Z(n117) );
  GTECH_OAI21 U113 ( .A(n126), .B(n127), .C(n128), .Z(n111) );
  GTECH_OAI21 U114 ( .A(n129), .B(n130), .C(n131), .Z(n128) );
  GTECH_NOT U115 ( .A(n130), .Z(n126) );
  GTECH_NOT U116 ( .A(n132), .Z(n112) );
  GTECH_NAND2 U117 ( .A(I_b[7]), .B(I_a[5]), .Z(n132) );
  GTECH_NOT U118 ( .A(n108), .Z(n110) );
  GTECH_NAND2 U119 ( .A(I_b[6]), .B(I_a[6]), .Z(n108) );
  GTECH_ADD_ABC U120 ( .A(n133), .B(n134), .C(n135), .COUT(n114) );
  GTECH_NOT U121 ( .A(n136), .Z(n135) );
  GTECH_XOR3 U122 ( .A(n137), .B(n138), .C(n139), .Z(n134) );
  GTECH_AND2 U123 ( .A(I_a[7]), .B(I_b[5]), .Z(n125) );
  GTECH_NOT U124 ( .A(n120), .Z(n118) );
  GTECH_OAI21 U125 ( .A(n139), .B(n140), .C(n141), .Z(n120) );
  GTECH_OAI21 U126 ( .A(n137), .B(n142), .C(n138), .Z(n141) );
  GTECH_NOT U127 ( .A(n140), .Z(n137) );
  GTECH_NOT U128 ( .A(n142), .Z(n139) );
  GTECH_ADD_ABC U129 ( .A(n143), .B(n144), .C(n145), .COUT(n124) );
  GTECH_NOT U130 ( .A(n146), .Z(n145) );
  GTECH_OA22 U131 ( .A(n147), .B(n148), .C(n149), .D(n150), .Z(n144) );
  GTECH_OA21 U132 ( .A(n151), .B(n152), .C(n153), .Z(n143) );
  GTECH_XOR3 U133 ( .A(n154), .B(n146), .C(n155), .Z(N151) );
  GTECH_OA21 U134 ( .A(n151), .B(n152), .C(n153), .Z(n155) );
  GTECH_OAI21 U135 ( .A(n156), .B(n157), .C(n158), .Z(n153) );
  GTECH_XOR3 U136 ( .A(n136), .B(n133), .C(n159), .Z(n146) );
  GTECH_XOR3 U137 ( .A(n138), .B(n142), .C(n140), .Z(n159) );
  GTECH_NAND2 U138 ( .A(I_a[7]), .B(I_b[4]), .Z(n140) );
  GTECH_OAI21 U139 ( .A(n160), .B(n161), .C(n162), .Z(n142) );
  GTECH_OAI21 U140 ( .A(n163), .B(n164), .C(n165), .Z(n162) );
  GTECH_NOT U141 ( .A(n166), .Z(n138) );
  GTECH_NAND2 U142 ( .A(I_a[6]), .B(I_b[5]), .Z(n166) );
  GTECH_ADD_ABC U143 ( .A(n167), .B(n168), .C(n169), .COUT(n133) );
  GTECH_NOT U144 ( .A(n170), .Z(n169) );
  GTECH_XOR3 U145 ( .A(n163), .B(n165), .C(n160), .Z(n168) );
  GTECH_NOT U146 ( .A(n164), .Z(n160) );
  GTECH_NOT U147 ( .A(n161), .Z(n163) );
  GTECH_XOR3 U148 ( .A(n129), .B(n131), .C(n130), .Z(n136) );
  GTECH_OAI21 U149 ( .A(n171), .B(n172), .C(n173), .Z(n130) );
  GTECH_OAI21 U150 ( .A(n174), .B(n175), .C(n176), .Z(n173) );
  GTECH_NOT U151 ( .A(n175), .Z(n171) );
  GTECH_NOT U152 ( .A(n177), .Z(n131) );
  GTECH_NAND2 U153 ( .A(I_b[7]), .B(I_a[4]), .Z(n177) );
  GTECH_NOT U154 ( .A(n127), .Z(n129) );
  GTECH_NAND2 U155 ( .A(I_b[6]), .B(I_a[5]), .Z(n127) );
  GTECH_OA22 U156 ( .A(n147), .B(n148), .C(n149), .D(n150), .Z(n154) );
  GTECH_NOT U157 ( .A(I_a[7]), .Z(n148) );
  GTECH_XOR3 U158 ( .A(n151), .B(n156), .C(n178), .Z(N150) );
  GTECH_NOT U159 ( .A(n158), .Z(n178) );
  GTECH_XOR3 U160 ( .A(n170), .B(n167), .C(n179), .Z(n158) );
  GTECH_XOR3 U161 ( .A(n165), .B(n164), .C(n161), .Z(n179) );
  GTECH_NAND2 U162 ( .A(I_a[6]), .B(I_b[4]), .Z(n161) );
  GTECH_OAI21 U163 ( .A(n180), .B(n181), .C(n182), .Z(n164) );
  GTECH_OAI21 U164 ( .A(n183), .B(n184), .C(n185), .Z(n182) );
  GTECH_NOT U165 ( .A(n186), .Z(n165) );
  GTECH_NAND2 U166 ( .A(I_a[5]), .B(I_b[5]), .Z(n186) );
  GTECH_ADD_ABC U167 ( .A(n187), .B(n188), .C(n189), .COUT(n167) );
  GTECH_NOT U168 ( .A(n190), .Z(n189) );
  GTECH_XOR3 U169 ( .A(n183), .B(n185), .C(n180), .Z(n188) );
  GTECH_NOT U170 ( .A(n184), .Z(n180) );
  GTECH_NOT U171 ( .A(n181), .Z(n183) );
  GTECH_XOR3 U172 ( .A(n174), .B(n176), .C(n175), .Z(n170) );
  GTECH_OAI21 U173 ( .A(n191), .B(n192), .C(n193), .Z(n175) );
  GTECH_OAI21 U174 ( .A(n194), .B(n195), .C(n196), .Z(n193) );
  GTECH_NOT U175 ( .A(n195), .Z(n191) );
  GTECH_NOT U176 ( .A(n197), .Z(n176) );
  GTECH_NAND2 U177 ( .A(I_b[7]), .B(I_a[3]), .Z(n197) );
  GTECH_NOT U178 ( .A(n172), .Z(n174) );
  GTECH_NAND2 U179 ( .A(I_b[6]), .B(I_a[4]), .Z(n172) );
  GTECH_NOT U180 ( .A(n152), .Z(n156) );
  GTECH_XNOR2 U181 ( .A(n149), .B(n150), .Z(n152) );
  GTECH_XNOR2 U182 ( .A(n147), .B(n198), .Z(n150) );
  GTECH_NAND2 U183 ( .A(I_a[7]), .B(I_b[3]), .Z(n198) );
  GTECH_AND2 U184 ( .A(n199), .B(n200), .Z(n147) );
  GTECH_OR_NOT U185 ( .A(n201), .B(n202), .Z(n200) );
  GTECH_OAI21 U186 ( .A(n203), .B(n202), .C(n204), .Z(n199) );
  GTECH_AOI2N2 U187 ( .A(n205), .B(n206), .C(n207), .D(n208), .Z(n149) );
  GTECH_NAND2 U188 ( .A(n207), .B(n208), .Z(n206) );
  GTECH_NOT U189 ( .A(n157), .Z(n151) );
  GTECH_OAI2N2 U190 ( .A(n209), .B(n210), .C(n211), .D(n212), .Z(n157) );
  GTECH_NAND2 U191 ( .A(n209), .B(n210), .Z(n212) );
  GTECH_XOR3 U192 ( .A(n209), .B(n213), .C(n214), .Z(N149) );
  GTECH_NOT U193 ( .A(n211), .Z(n214) );
  GTECH_XOR3 U194 ( .A(n190), .B(n187), .C(n215), .Z(n211) );
  GTECH_XOR3 U195 ( .A(n185), .B(n184), .C(n181), .Z(n215) );
  GTECH_NAND2 U196 ( .A(I_a[5]), .B(I_b[4]), .Z(n181) );
  GTECH_OAI21 U197 ( .A(n216), .B(n217), .C(n218), .Z(n184) );
  GTECH_OAI21 U198 ( .A(n219), .B(n220), .C(n221), .Z(n218) );
  GTECH_NOT U199 ( .A(n222), .Z(n185) );
  GTECH_NAND2 U200 ( .A(I_b[5]), .B(I_a[4]), .Z(n222) );
  GTECH_ADD_ABC U201 ( .A(n223), .B(n224), .C(n225), .COUT(n187) );
  GTECH_XOR3 U202 ( .A(n219), .B(n221), .C(n216), .Z(n224) );
  GTECH_NOT U203 ( .A(n220), .Z(n216) );
  GTECH_OA21 U204 ( .A(n226), .B(n227), .C(n228), .Z(n223) );
  GTECH_XOR3 U205 ( .A(n194), .B(n196), .C(n195), .Z(n190) );
  GTECH_OAI21 U206 ( .A(n229), .B(n230), .C(n231), .Z(n195) );
  GTECH_NOT U207 ( .A(n232), .Z(n196) );
  GTECH_NAND2 U208 ( .A(I_b[7]), .B(I_a[2]), .Z(n232) );
  GTECH_NOT U209 ( .A(n192), .Z(n194) );
  GTECH_NAND2 U210 ( .A(I_b[6]), .B(I_a[3]), .Z(n192) );
  GTECH_NOT U211 ( .A(n210), .Z(n213) );
  GTECH_XOR3 U212 ( .A(n233), .B(n207), .C(n205), .Z(n210) );
  GTECH_XOR3 U213 ( .A(n203), .B(n204), .C(n202), .Z(n205) );
  GTECH_OAI21 U214 ( .A(n234), .B(n235), .C(n236), .Z(n202) );
  GTECH_OAI21 U215 ( .A(n237), .B(n238), .C(n239), .Z(n236) );
  GTECH_NOT U216 ( .A(n238), .Z(n234) );
  GTECH_NOT U217 ( .A(n240), .Z(n204) );
  GTECH_NAND2 U218 ( .A(I_a[6]), .B(I_b[3]), .Z(n240) );
  GTECH_NOT U219 ( .A(n201), .Z(n203) );
  GTECH_NAND2 U220 ( .A(I_a[7]), .B(I_b[2]), .Z(n201) );
  GTECH_ADD_ABC U221 ( .A(n241), .B(n242), .C(n243), .COUT(n207) );
  GTECH_XNOR2 U222 ( .A(n244), .B(n245), .Z(n242) );
  GTECH_NAND2 U223 ( .A(I_a[7]), .B(I_b[1]), .Z(n245) );
  GTECH_NOT U224 ( .A(n208), .Z(n233) );
  GTECH_NAND2 U225 ( .A(I_a[7]), .B(n246), .Z(n208) );
  GTECH_ADD_ABC U226 ( .A(n247), .B(n248), .C(n249), .COUT(n209) );
  GTECH_XOR3 U227 ( .A(n241), .B(n250), .C(n243), .Z(n248) );
  GTECH_NOT U228 ( .A(n251), .Z(n243) );
  GTECH_XOR3 U229 ( .A(n252), .B(n249), .C(n247), .Z(N148) );
  GTECH_ADD_ABC U230 ( .A(n253), .B(n254), .C(n255), .COUT(n247) );
  GTECH_NOT U231 ( .A(n256), .Z(n255) );
  GTECH_XOR3 U232 ( .A(n257), .B(n258), .C(n259), .Z(n254) );
  GTECH_NOT U233 ( .A(n260), .Z(n258) );
  GTECH_XOR3 U234 ( .A(n261), .B(n225), .C(n262), .Z(n249) );
  GTECH_OAI21 U235 ( .A(n226), .B(n227), .C(n228), .Z(n262) );
  GTECH_OAI21 U236 ( .A(n263), .B(n264), .C(n265), .Z(n228) );
  GTECH_NOT U237 ( .A(n226), .Z(n264) );
  GTECH_XOR3 U238 ( .A(n266), .B(n267), .C(n231), .Z(n225) );
  GTECH_NAND3 U239 ( .A(I_b[6]), .B(I_a[1]), .C(n268), .Z(n231) );
  GTECH_NOT U240 ( .A(n230), .Z(n267) );
  GTECH_NAND2 U241 ( .A(I_b[7]), .B(I_a[1]), .Z(n230) );
  GTECH_NOT U242 ( .A(n229), .Z(n266) );
  GTECH_NAND2 U243 ( .A(I_b[6]), .B(I_a[2]), .Z(n229) );
  GTECH_XOR3 U244 ( .A(n221), .B(n220), .C(n219), .Z(n261) );
  GTECH_NOT U245 ( .A(n217), .Z(n219) );
  GTECH_NAND2 U246 ( .A(I_b[4]), .B(I_a[4]), .Z(n217) );
  GTECH_OAI21 U247 ( .A(n269), .B(n270), .C(n271), .Z(n220) );
  GTECH_OAI21 U248 ( .A(n272), .B(n273), .C(n274), .Z(n271) );
  GTECH_NOT U249 ( .A(n273), .Z(n269) );
  GTECH_NOT U250 ( .A(n275), .Z(n221) );
  GTECH_NAND2 U251 ( .A(I_b[5]), .B(I_a[3]), .Z(n275) );
  GTECH_XOR3 U252 ( .A(n250), .B(n251), .C(n241), .Z(n252) );
  GTECH_ADD_ABC U253 ( .A(n257), .B(n276), .C(n259), .COUT(n241) );
  GTECH_NOT U254 ( .A(n277), .Z(n259) );
  GTECH_XOR3 U255 ( .A(n278), .B(n279), .C(n280), .Z(n276) );
  GTECH_XOR3 U256 ( .A(n237), .B(n239), .C(n238), .Z(n251) );
  GTECH_OAI21 U257 ( .A(n281), .B(n282), .C(n283), .Z(n238) );
  GTECH_OAI21 U258 ( .A(n284), .B(n285), .C(n286), .Z(n283) );
  GTECH_NOT U259 ( .A(n285), .Z(n281) );
  GTECH_NOT U260 ( .A(n287), .Z(n239) );
  GTECH_NAND2 U261 ( .A(I_a[5]), .B(I_b[3]), .Z(n287) );
  GTECH_NOT U262 ( .A(n235), .Z(n237) );
  GTECH_NAND2 U263 ( .A(I_a[6]), .B(I_b[2]), .Z(n235) );
  GTECH_XNOR2 U264 ( .A(n244), .B(n288), .Z(n250) );
  GTECH_NAND2 U265 ( .A(I_a[7]), .B(I_b[1]), .Z(n288) );
  GTECH_NOT U266 ( .A(n246), .Z(n244) );
  GTECH_OAI21 U267 ( .A(n280), .B(n289), .C(n290), .Z(n246) );
  GTECH_OAI21 U268 ( .A(n278), .B(n291), .C(n279), .Z(n290) );
  GTECH_NOT U269 ( .A(n291), .Z(n280) );
  GTECH_XOR3 U270 ( .A(n256), .B(n253), .C(n292), .Z(N147) );
  GTECH_XOR3 U271 ( .A(n277), .B(n257), .C(n260), .Z(n292) );
  GTECH_XOR3 U272 ( .A(n278), .B(n279), .C(n291), .Z(n260) );
  GTECH_OAI21 U273 ( .A(n293), .B(n294), .C(n295), .Z(n291) );
  GTECH_OAI21 U274 ( .A(n296), .B(n297), .C(n298), .Z(n295) );
  GTECH_NOT U275 ( .A(n299), .Z(n279) );
  GTECH_NAND2 U276 ( .A(I_a[6]), .B(I_b[1]), .Z(n299) );
  GTECH_NOT U277 ( .A(n289), .Z(n278) );
  GTECH_NAND2 U278 ( .A(I_a[7]), .B(I_b[0]), .Z(n289) );
  GTECH_ADD_ABC U279 ( .A(n300), .B(n301), .C(n302), .COUT(n257) );
  GTECH_XOR3 U280 ( .A(n296), .B(n298), .C(n293), .Z(n301) );
  GTECH_NOT U281 ( .A(n297), .Z(n293) );
  GTECH_XOR3 U282 ( .A(n284), .B(n286), .C(n285), .Z(n277) );
  GTECH_OAI21 U283 ( .A(n303), .B(n304), .C(n305), .Z(n285) );
  GTECH_OAI21 U284 ( .A(n306), .B(n307), .C(n308), .Z(n305) );
  GTECH_NOT U285 ( .A(n307), .Z(n303) );
  GTECH_NOT U286 ( .A(n309), .Z(n286) );
  GTECH_NAND2 U287 ( .A(I_b[3]), .B(I_a[4]), .Z(n309) );
  GTECH_NOT U288 ( .A(n282), .Z(n284) );
  GTECH_NAND2 U289 ( .A(I_a[5]), .B(I_b[2]), .Z(n282) );
  GTECH_ADD_ABC U290 ( .A(n310), .B(n311), .C(n312), .COUT(n253) );
  GTECH_XOR3 U291 ( .A(n300), .B(n313), .C(n302), .Z(n311) );
  GTECH_NOT U292 ( .A(n314), .Z(n302) );
  GTECH_OA21 U293 ( .A(n315), .B(n316), .C(n317), .Z(n310) );
  GTECH_XOR3 U294 ( .A(n265), .B(n227), .C(n226), .Z(n256) );
  GTECH_XNOR2 U295 ( .A(n268), .B(n318), .Z(n226) );
  GTECH_AND2 U296 ( .A(I_b[6]), .B(I_a[1]), .Z(n318) );
  GTECH_NOT U297 ( .A(n319), .Z(n268) );
  GTECH_NAND2 U298 ( .A(I_b[7]), .B(I_a[0]), .Z(n319) );
  GTECH_NOT U299 ( .A(n263), .Z(n227) );
  GTECH_XOR3 U300 ( .A(n272), .B(n274), .C(n273), .Z(n263) );
  GTECH_OAI21 U301 ( .A(n320), .B(n321), .C(n322), .Z(n273) );
  GTECH_NOT U302 ( .A(n323), .Z(n274) );
  GTECH_NAND2 U303 ( .A(I_b[5]), .B(I_a[2]), .Z(n323) );
  GTECH_NOT U304 ( .A(n270), .Z(n272) );
  GTECH_NAND2 U305 ( .A(I_b[4]), .B(I_a[3]), .Z(n270) );
  GTECH_NOT U306 ( .A(n324), .Z(n265) );
  GTECH_NAND3 U307 ( .A(I_a[0]), .B(n325), .C(I_b[6]), .Z(n324) );
  GTECH_XOR3 U308 ( .A(n326), .B(n312), .C(n327), .Z(N146) );
  GTECH_OA21 U309 ( .A(n315), .B(n316), .C(n317), .Z(n327) );
  GTECH_OAI21 U310 ( .A(n328), .B(n329), .C(n330), .Z(n317) );
  GTECH_NOT U311 ( .A(n315), .Z(n329) );
  GTECH_XNOR2 U312 ( .A(n331), .B(n325), .Z(n312) );
  GTECH_NOT U313 ( .A(n332), .Z(n325) );
  GTECH_XOR3 U314 ( .A(n333), .B(n334), .C(n322), .Z(n332) );
  GTECH_NAND3 U315 ( .A(I_b[4]), .B(I_a[1]), .C(n335), .Z(n322) );
  GTECH_NOT U316 ( .A(n321), .Z(n334) );
  GTECH_NAND2 U317 ( .A(I_b[5]), .B(I_a[1]), .Z(n321) );
  GTECH_NOT U318 ( .A(n320), .Z(n333) );
  GTECH_NAND2 U319 ( .A(I_b[4]), .B(I_a[2]), .Z(n320) );
  GTECH_AND2 U320 ( .A(I_b[6]), .B(I_a[0]), .Z(n331) );
  GTECH_XOR3 U321 ( .A(n313), .B(n314), .C(n300), .Z(n326) );
  GTECH_ADD_ABC U322 ( .A(n336), .B(n337), .C(n338), .COUT(n300) );
  GTECH_NOT U323 ( .A(n339), .Z(n338) );
  GTECH_XOR3 U324 ( .A(n340), .B(n341), .C(n342), .Z(n337) );
  GTECH_XOR3 U325 ( .A(n306), .B(n308), .C(n307), .Z(n314) );
  GTECH_OAI21 U326 ( .A(n343), .B(n344), .C(n345), .Z(n307) );
  GTECH_OAI21 U327 ( .A(n346), .B(n347), .C(n348), .Z(n345) );
  GTECH_NOT U328 ( .A(n347), .Z(n343) );
  GTECH_NOT U329 ( .A(n349), .Z(n308) );
  GTECH_NAND2 U330 ( .A(I_b[3]), .B(I_a[3]), .Z(n349) );
  GTECH_NOT U331 ( .A(n304), .Z(n306) );
  GTECH_NAND2 U332 ( .A(I_b[2]), .B(I_a[4]), .Z(n304) );
  GTECH_NOT U333 ( .A(n350), .Z(n313) );
  GTECH_XOR3 U334 ( .A(n296), .B(n298), .C(n297), .Z(n350) );
  GTECH_OAI21 U335 ( .A(n342), .B(n351), .C(n352), .Z(n297) );
  GTECH_OAI21 U336 ( .A(n340), .B(n353), .C(n341), .Z(n352) );
  GTECH_NOT U337 ( .A(n351), .Z(n340) );
  GTECH_NOT U338 ( .A(n353), .Z(n342) );
  GTECH_NOT U339 ( .A(n354), .Z(n298) );
  GTECH_NAND2 U340 ( .A(I_a[5]), .B(I_b[1]), .Z(n354) );
  GTECH_NOT U341 ( .A(n294), .Z(n296) );
  GTECH_NAND2 U342 ( .A(I_a[6]), .B(I_b[0]), .Z(n294) );
  GTECH_XOR3 U343 ( .A(n330), .B(n316), .C(n315), .Z(N145) );
  GTECH_XNOR2 U344 ( .A(n335), .B(n355), .Z(n315) );
  GTECH_AND2 U345 ( .A(I_b[4]), .B(I_a[1]), .Z(n355) );
  GTECH_NOT U346 ( .A(n356), .Z(n335) );
  GTECH_NAND2 U347 ( .A(I_b[5]), .B(I_a[0]), .Z(n356) );
  GTECH_NOT U348 ( .A(n328), .Z(n316) );
  GTECH_XOR3 U349 ( .A(n339), .B(n336), .C(n357), .Z(n328) );
  GTECH_XOR3 U350 ( .A(n341), .B(n353), .C(n351), .Z(n357) );
  GTECH_NAND2 U351 ( .A(I_a[5]), .B(I_b[0]), .Z(n351) );
  GTECH_OAI21 U352 ( .A(n358), .B(n359), .C(n360), .Z(n353) );
  GTECH_OAI21 U353 ( .A(n361), .B(n362), .C(n363), .Z(n360) );
  GTECH_NOT U354 ( .A(n364), .Z(n341) );
  GTECH_NAND2 U355 ( .A(I_a[4]), .B(I_b[1]), .Z(n364) );
  GTECH_ADD_ABC U356 ( .A(n365), .B(n366), .C(n367), .COUT(n336) );
  GTECH_XOR3 U357 ( .A(n361), .B(n363), .C(n358), .Z(n366) );
  GTECH_NOT U358 ( .A(n362), .Z(n358) );
  GTECH_OA21 U359 ( .A(n368), .B(n369), .C(n370), .Z(n365) );
  GTECH_XOR3 U360 ( .A(n346), .B(n348), .C(n347), .Z(n339) );
  GTECH_OAI21 U361 ( .A(n371), .B(n372), .C(n373), .Z(n347) );
  GTECH_NOT U362 ( .A(n374), .Z(n348) );
  GTECH_NAND2 U363 ( .A(I_b[3]), .B(I_a[2]), .Z(n374) );
  GTECH_NOT U364 ( .A(n344), .Z(n346) );
  GTECH_NAND2 U365 ( .A(I_b[2]), .B(I_a[3]), .Z(n344) );
  GTECH_NOT U366 ( .A(n375), .Z(n330) );
  GTECH_NAND3 U367 ( .A(I_a[0]), .B(n376), .C(I_b[4]), .Z(n375) );
  GTECH_NOT U368 ( .A(n377), .Z(n376) );
  GTECH_XNOR2 U369 ( .A(n378), .B(n377), .Z(N144) );
  GTECH_XOR3 U370 ( .A(n379), .B(n367), .C(n380), .Z(n377) );
  GTECH_OAI21 U371 ( .A(n368), .B(n369), .C(n370), .Z(n380) );
  GTECH_OAI21 U372 ( .A(n381), .B(n382), .C(n383), .Z(n370) );
  GTECH_NOT U373 ( .A(n368), .Z(n382) );
  GTECH_XOR3 U374 ( .A(n384), .B(n385), .C(n373), .Z(n367) );
  GTECH_NAND3 U375 ( .A(I_b[2]), .B(I_a[1]), .C(n386), .Z(n373) );
  GTECH_NOT U376 ( .A(n372), .Z(n385) );
  GTECH_NAND2 U377 ( .A(I_b[3]), .B(I_a[1]), .Z(n372) );
  GTECH_NOT U378 ( .A(n371), .Z(n384) );
  GTECH_NAND2 U379 ( .A(I_b[2]), .B(I_a[2]), .Z(n371) );
  GTECH_XOR3 U380 ( .A(n363), .B(n362), .C(n361), .Z(n379) );
  GTECH_NOT U381 ( .A(n359), .Z(n361) );
  GTECH_NAND2 U382 ( .A(I_a[4]), .B(I_b[0]), .Z(n359) );
  GTECH_OAI21 U383 ( .A(n387), .B(n388), .C(n389), .Z(n362) );
  GTECH_OAI21 U384 ( .A(n390), .B(n391), .C(n392), .Z(n389) );
  GTECH_NOT U385 ( .A(n391), .Z(n387) );
  GTECH_NOT U386 ( .A(n393), .Z(n363) );
  GTECH_NAND2 U387 ( .A(I_a[3]), .B(I_b[1]), .Z(n393) );
  GTECH_AND2 U388 ( .A(I_b[4]), .B(I_a[0]), .Z(n378) );
  GTECH_XOR3 U389 ( .A(n383), .B(n369), .C(n368), .Z(N143) );
  GTECH_XNOR2 U390 ( .A(n386), .B(n394), .Z(n368) );
  GTECH_AND2 U391 ( .A(I_b[2]), .B(I_a[1]), .Z(n394) );
  GTECH_NOT U392 ( .A(n395), .Z(n386) );
  GTECH_NAND2 U393 ( .A(I_b[3]), .B(I_a[0]), .Z(n395) );
  GTECH_NOT U394 ( .A(n381), .Z(n369) );
  GTECH_XOR3 U395 ( .A(n390), .B(n392), .C(n391), .Z(n381) );
  GTECH_OAI21 U396 ( .A(n396), .B(n397), .C(n398), .Z(n391) );
  GTECH_NOT U397 ( .A(n399), .Z(n392) );
  GTECH_NAND2 U398 ( .A(I_b[1]), .B(I_a[2]), .Z(n399) );
  GTECH_NOT U399 ( .A(n388), .Z(n390) );
  GTECH_NAND2 U400 ( .A(I_b[0]), .B(I_a[3]), .Z(n388) );
  GTECH_NOT U401 ( .A(n400), .Z(n383) );
  GTECH_NAND3 U402 ( .A(I_a[0]), .B(n401), .C(I_b[2]), .Z(n400) );
  GTECH_NOT U403 ( .A(n402), .Z(n401) );
  GTECH_XNOR2 U404 ( .A(n403), .B(n402), .Z(N142) );
  GTECH_XOR3 U405 ( .A(n404), .B(n405), .C(n398), .Z(n402) );
  GTECH_NAND3 U406 ( .A(n406), .B(I_b[0]), .C(I_a[1]), .Z(n398) );
  GTECH_NOT U407 ( .A(n396), .Z(n405) );
  GTECH_NAND2 U408 ( .A(I_a[1]), .B(I_b[1]), .Z(n396) );
  GTECH_NOT U409 ( .A(n397), .Z(n404) );
  GTECH_NAND2 U410 ( .A(I_b[0]), .B(I_a[2]), .Z(n397) );
  GTECH_AND2 U411 ( .A(I_b[2]), .B(I_a[0]), .Z(n403) );
  GTECH_XNOR2 U412 ( .A(n406), .B(n407), .Z(N141) );
  GTECH_NAND2 U413 ( .A(I_a[1]), .B(I_b[0]), .Z(n407) );
  GTECH_NOT U414 ( .A(n408), .Z(n406) );
  GTECH_NAND2 U415 ( .A(I_a[0]), .B(I_b[1]), .Z(n408) );
  GTECH_AND2 U416 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

