
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374;

  GTECH_MUX2 U137 ( .A(n276), .B(n277), .S(n278), .Z(sum[9]) );
  GTECH_OA21 U138 ( .A(n279), .B(n280), .C(n281), .Z(n278) );
  GTECH_ADD_AB U139 ( .A(b[9]), .B(a[9]), .S(n277) );
  GTECH_OR_NOT U140 ( .A(n282), .B(n283), .Z(n276) );
  GTECH_NAND2 U141 ( .A(n284), .B(n285), .Z(sum[8]) );
  GTECH_AO21 U142 ( .A(n281), .B(n286), .C(n280), .Z(n284) );
  GTECH_MUX2 U143 ( .A(n287), .B(n288), .S(n289), .Z(sum[7]) );
  GTECH_ADD_AB U144 ( .A(n290), .B(n291), .S(n288) );
  GTECH_XNOR2 U145 ( .A(n292), .B(n291), .Z(n287) );
  GTECH_ADD_AB U146 ( .A(b[7]), .B(a[7]), .S(n291) );
  GTECH_OA21 U147 ( .A(n293), .B(n294), .C(n295), .Z(n292) );
  GTECH_MUX2 U148 ( .A(n296), .B(n297), .S(n289), .Z(sum[6]) );
  GTECH_XNOR2 U149 ( .A(n298), .B(n299), .Z(n297) );
  GTECH_XNOR2 U150 ( .A(n294), .B(n299), .Z(n296) );
  GTECH_AND2 U151 ( .A(n295), .B(n300), .Z(n299) );
  GTECH_AOI21 U152 ( .A(n301), .B(n302), .C(n303), .Z(n294) );
  GTECH_XNOR2 U153 ( .A(n304), .B(n305), .Z(sum[5]) );
  GTECH_OR_NOT U154 ( .A(n303), .B(n301), .Z(n305) );
  GTECH_OA21 U155 ( .A(n302), .B(n289), .C(n306), .Z(n304) );
  GTECH_XNOR2 U156 ( .A(n307), .B(n289), .Z(sum[4]) );
  GTECH_MUX2 U157 ( .A(n308), .B(n309), .S(cin), .Z(sum[3]) );
  GTECH_ADD_AB U158 ( .A(n310), .B(n311), .S(n309) );
  GTECH_XNOR2 U159 ( .A(n312), .B(n311), .Z(n308) );
  GTECH_ADD_AB U160 ( .A(b[3]), .B(a[3]), .S(n311) );
  GTECH_OA21 U161 ( .A(n313), .B(n314), .C(n315), .Z(n312) );
  GTECH_MUX2 U162 ( .A(n316), .B(n317), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U163 ( .A(n318), .B(n319), .Z(n317) );
  GTECH_XNOR2 U164 ( .A(n319), .B(n314), .Z(n316) );
  GTECH_AOI21 U165 ( .A(n320), .B(n321), .C(n322), .Z(n314) );
  GTECH_AND2 U166 ( .A(n315), .B(n323), .Z(n319) );
  GTECH_MUX2 U167 ( .A(n324), .B(n325), .S(n326), .Z(sum[1]) );
  GTECH_AND_NOT U168 ( .A(n320), .B(n322), .Z(n326) );
  GTECH_OAI21 U169 ( .A(cin), .B(n321), .C(n327), .Z(n325) );
  GTECH_AO21 U170 ( .A(n327), .B(cin), .C(n321), .Z(n324) );
  GTECH_MUX2 U171 ( .A(n328), .B(n329), .S(n330), .Z(sum[15]) );
  GTECH_ADD_AB U172 ( .A(n331), .B(n332), .S(n329) );
  GTECH_XNOR2 U173 ( .A(n333), .B(n332), .Z(n328) );
  GTECH_ADD_AB U174 ( .A(b[15]), .B(a[15]), .S(n332) );
  GTECH_OA21 U175 ( .A(n334), .B(n335), .C(n336), .Z(n333) );
  GTECH_MUX2 U176 ( .A(n337), .B(n338), .S(n330), .Z(sum[14]) );
  GTECH_XNOR2 U177 ( .A(n339), .B(n340), .Z(n338) );
  GTECH_XNOR2 U178 ( .A(n340), .B(n335), .Z(n337) );
  GTECH_AOI21 U179 ( .A(n341), .B(n342), .C(n343), .Z(n335) );
  GTECH_AND2 U180 ( .A(n336), .B(n344), .Z(n340) );
  GTECH_MUX2 U181 ( .A(n345), .B(n346), .S(n347), .Z(sum[13]) );
  GTECH_AOI21 U182 ( .A(n330), .B(n348), .C(n342), .Z(n347) );
  GTECH_NOT U183 ( .A(n349), .Z(n330) );
  GTECH_ADD_AB U184 ( .A(b[13]), .B(a[13]), .S(n346) );
  GTECH_OR_NOT U185 ( .A(n343), .B(n341), .Z(n345) );
  GTECH_NAND2 U186 ( .A(n350), .B(n351), .Z(sum[12]) );
  GTECH_AO21 U187 ( .A(n352), .B(n348), .C(n349), .Z(n350) );
  GTECH_MUX2 U188 ( .A(n353), .B(n354), .S(n280), .Z(sum[11]) );
  GTECH_XNOR2 U189 ( .A(n355), .B(n356), .Z(n354) );
  GTECH_OA21 U190 ( .A(a[10]), .B(n357), .C(n358), .Z(n355) );
  GTECH_AO21 U191 ( .A(n357), .B(a[10]), .C(b[10]), .Z(n358) );
  GTECH_XNOR2 U192 ( .A(n359), .B(n356), .Z(n353) );
  GTECH_XNOR2 U193 ( .A(b[11]), .B(a[11]), .Z(n356) );
  GTECH_MUX2 U194 ( .A(n360), .B(n361), .S(n280), .Z(sum[10]) );
  GTECH_ADD_AB U195 ( .A(n357), .B(n362), .S(n361) );
  GTECH_OAI21 U196 ( .A(n282), .B(n281), .C(n283), .Z(n357) );
  GTECH_ADD_AB U197 ( .A(n363), .B(n362), .S(n360) );
  GTECH_ADD_AB U198 ( .A(b[10]), .B(a[10]), .S(n362) );
  GTECH_ADD_AB U199 ( .A(cin), .B(n364), .S(sum[0]) );
  GTECH_OAI21 U200 ( .A(n349), .B(n365), .C(n351), .Z(cout) );
  GTECH_NAND3 U201 ( .A(n348), .B(n352), .C(n349), .Z(n351) );
  GTECH_NOT U202 ( .A(n342), .Z(n352) );
  GTECH_AND2 U203 ( .A(a[12]), .B(b[12]), .Z(n342) );
  GTECH_AOI21 U204 ( .A(n331), .B(a[15]), .C(n366), .Z(n365) );
  GTECH_OA21 U205 ( .A(a[15]), .B(n331), .C(b[15]), .Z(n366) );
  GTECH_OAI21 U206 ( .A(n339), .B(n334), .C(n336), .Z(n331) );
  GTECH_NAND2 U207 ( .A(a[14]), .B(b[14]), .Z(n336) );
  GTECH_NOT U208 ( .A(n344), .Z(n334) );
  GTECH_OR2 U209 ( .A(a[14]), .B(b[14]), .Z(n344) );
  GTECH_AOI21 U210 ( .A(n341), .B(n348), .C(n343), .Z(n339) );
  GTECH_AND2 U211 ( .A(b[13]), .B(a[13]), .Z(n343) );
  GTECH_OR2 U212 ( .A(a[12]), .B(b[12]), .Z(n348) );
  GTECH_OR2 U213 ( .A(b[13]), .B(a[13]), .Z(n341) );
  GTECH_OA21 U214 ( .A(n367), .B(n280), .C(n285), .Z(n349) );
  GTECH_NAND3 U215 ( .A(n286), .B(n281), .C(n280), .Z(n285) );
  GTECH_NAND2 U216 ( .A(b[8]), .B(a[8]), .Z(n281) );
  GTECH_MUX2 U217 ( .A(n307), .B(n368), .S(n289), .Z(n280) );
  GTECH_MUX2 U218 ( .A(n364), .B(n369), .S(cin), .Z(n289) );
  GTECH_OA21 U219 ( .A(a[3]), .B(n310), .C(n370), .Z(n369) );
  GTECH_AO21 U220 ( .A(n310), .B(a[3]), .C(b[3]), .Z(n370) );
  GTECH_OAI21 U221 ( .A(n318), .B(n313), .C(n315), .Z(n310) );
  GTECH_NAND2 U222 ( .A(a[2]), .B(b[2]), .Z(n315) );
  GTECH_NOT U223 ( .A(n323), .Z(n313) );
  GTECH_OR2 U224 ( .A(a[2]), .B(b[2]), .Z(n323) );
  GTECH_AOI21 U225 ( .A(n320), .B(n327), .C(n322), .Z(n318) );
  GTECH_AND2 U226 ( .A(b[1]), .B(a[1]), .Z(n322) );
  GTECH_OR2 U227 ( .A(b[1]), .B(a[1]), .Z(n320) );
  GTECH_AND_NOT U228 ( .A(n327), .B(n321), .Z(n364) );
  GTECH_AND2 U229 ( .A(b[0]), .B(a[0]), .Z(n321) );
  GTECH_OR2 U230 ( .A(a[0]), .B(b[0]), .Z(n327) );
  GTECH_AOI21 U231 ( .A(n290), .B(a[7]), .C(n371), .Z(n368) );
  GTECH_OA21 U232 ( .A(a[7]), .B(n290), .C(b[7]), .Z(n371) );
  GTECH_OAI21 U233 ( .A(n298), .B(n293), .C(n295), .Z(n290) );
  GTECH_NAND2 U234 ( .A(a[6]), .B(b[6]), .Z(n295) );
  GTECH_NOT U235 ( .A(n300), .Z(n293) );
  GTECH_OR2 U236 ( .A(a[6]), .B(b[6]), .Z(n300) );
  GTECH_AOI21 U237 ( .A(n306), .B(n301), .C(n303), .Z(n298) );
  GTECH_AND2 U238 ( .A(b[5]), .B(a[5]), .Z(n303) );
  GTECH_OR2 U239 ( .A(a[5]), .B(b[5]), .Z(n301) );
  GTECH_OR_NOT U240 ( .A(n302), .B(n306), .Z(n307) );
  GTECH_OR2 U241 ( .A(b[4]), .B(a[4]), .Z(n306) );
  GTECH_AND2 U242 ( .A(a[4]), .B(b[4]), .Z(n302) );
  GTECH_AOI21 U243 ( .A(n359), .B(a[11]), .C(n372), .Z(n367) );
  GTECH_OA21 U244 ( .A(a[11]), .B(n359), .C(b[11]), .Z(n372) );
  GTECH_AO21 U245 ( .A(n363), .B(a[10]), .C(n373), .Z(n359) );
  GTECH_OA21 U246 ( .A(a[10]), .B(n363), .C(b[10]), .Z(n373) );
  GTECH_OAI21 U247 ( .A(n282), .B(n279), .C(n283), .Z(n363) );
  GTECH_OR_NOT U248 ( .A(n374), .B(b[9]), .Z(n283) );
  GTECH_NOT U249 ( .A(n286), .Z(n279) );
  GTECH_OR2 U250 ( .A(a[8]), .B(b[8]), .Z(n286) );
  GTECH_AND_NOT U251 ( .A(n374), .B(b[9]), .Z(n282) );
  GTECH_NOT U252 ( .A(a[9]), .Z(n374) );
endmodule

