
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n117, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n117), .K(n117), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n254) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n117), .K(n117), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n117), .K(n117), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n117), .K(n117), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n117), .K(n117), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n117), .K(n117), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]) );
  GTECH_FJK1S A_reg_15_ ( .J(n117), .K(n117), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n270) );
  GTECH_FJK1S A_reg_14_ ( .J(n117), .K(n117), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n269) );
  GTECH_FJK1S A_reg_13_ ( .J(n117), .K(n117), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n268) );
  GTECH_FJK1S A_reg_12_ ( .J(n117), .K(n117), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n267) );
  GTECH_FJK1S A_reg_11_ ( .J(n117), .K(n117), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n266) );
  GTECH_FJK1S A_reg_10_ ( .J(n117), .K(n117), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n265) );
  GTECH_FJK1S A_reg_9_ ( .J(n117), .K(n117), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n264) );
  GTECH_FJK1S A_reg_8_ ( .J(n117), .K(n117), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n263) );
  GTECH_FJK1S A_reg_7_ ( .J(n117), .K(n117), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n262) );
  GTECH_FJK1S A_reg_6_ ( .J(n117), .K(n117), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n261) );
  GTECH_FJK1S A_reg_5_ ( .J(n117), .K(n117), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n260) );
  GTECH_FJK1S A_reg_4_ ( .J(n117), .K(n117), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n259) );
  GTECH_FJK1S A_reg_3_ ( .J(n117), .K(n117), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n258) );
  GTECH_FJK1S A_reg_2_ ( .J(n117), .K(n117), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n257) );
  GTECH_FJK1S A_reg_1_ ( .J(n117), .K(n117), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n256) );
  GTECH_FJK1S A_reg_0_ ( .J(n117), .K(n117), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n255) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n117), .K(n117), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n117), .K(n117), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n117), .K(n117), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n117), .K(n117), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n117), .K(n117), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n117), .K(n117), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n117), .K(n117), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n117), .K(n117), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n117), .K(n117), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n117), .K(n117), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n117), .K(n117), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n117), .K(n117), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n117), .K(n117), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n117), .K(n117), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n117), .K(n117), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n117), .K(n117), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n117), .K(n117), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n117), .K(n117), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n117), .K(n117), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n117), .K(n117), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n117), .K(n117), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n117), .K(n117), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n117), .K(n117), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n117), .K(n117), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n117), .K(n117), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n117), .K(n117), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n117), .K(n117), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n117), .K(n117), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n117), .K(n117), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n117), .K(n117), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n117), .K(n117), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n117), .K(n117), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n117), .K(n117), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n117), .K(n117), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n117), .K(n117), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n117), .K(n117), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n117), .K(n117), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n117), .K(n117), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n117), .K(n117), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n117), .K(n117), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n117), .K(n117), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n117), .K(n117), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n117), .K(n117), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n117), .K(n117), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n117), .K(n117), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n117), .K(n117), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n117), .K(n117), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n117), .K(n117), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n117), .K(n117), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n117), .K(n117), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n117), .K(n117), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n117), .K(n117), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n117), .K(n117), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n117), .K(n117), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n117), .K(n117), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n117), .K(n117), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n117), .K(n117), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n117), .K(n117), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n117), .K(n117), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n117), .K(n117), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n117), .K(n117), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n117), .K(n117), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n117), .K(n117), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n117), .K(n117), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n117), .K(n117), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n117), .K(n117), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U256 ( .Z(n117) );
  GTECH_NOT U257 ( .A(n272), .Z(N99) );
  GTECH_AOI222 U258 ( .A(n273), .B(n274), .C(n275), .D(n276), .E(n277), .F(
        n278), .Z(n272) );
  GTECH_NOT U259 ( .A(n279), .Z(N98) );
  GTECH_AOI222 U260 ( .A(n273), .B(n280), .C(n281), .D(n282), .E(R[15]), .F(
        n283), .Z(n279) );
  GTECH_OR_NOT U261 ( .A(n275), .B(n284), .Z(n281) );
  GTECH_OAI2N2 U262 ( .A(n13), .B(n285), .C(R[14]), .D(n283), .Z(N97) );
  GTECH_OAI2N2 U263 ( .A(n14), .B(n285), .C(R[13]), .D(n283), .Z(N96) );
  GTECH_OAI2N2 U264 ( .A(n15), .B(n285), .C(R[12]), .D(n283), .Z(N95) );
  GTECH_OAI2N2 U265 ( .A(n16), .B(n285), .C(R[11]), .D(n283), .Z(N94) );
  GTECH_OAI2N2 U266 ( .A(n17), .B(n285), .C(R[10]), .D(n283), .Z(N93) );
  GTECH_OAI2N2 U267 ( .A(n18), .B(n285), .C(R[9]), .D(n283), .Z(N92) );
  GTECH_OAI2N2 U268 ( .A(n19), .B(n285), .C(R[8]), .D(n283), .Z(N91) );
  GTECH_OAI2N2 U269 ( .A(n20), .B(n285), .C(R[7]), .D(n283), .Z(N90) );
  GTECH_OAI2N2 U270 ( .A(n21), .B(n285), .C(R[6]), .D(n283), .Z(N89) );
  GTECH_OAI2N2 U271 ( .A(n22), .B(n285), .C(R[5]), .D(n283), .Z(N88) );
  GTECH_OAI2N2 U272 ( .A(n23), .B(n285), .C(R[4]), .D(n283), .Z(N87) );
  GTECH_OAI2N2 U273 ( .A(n24), .B(n285), .C(R[3]), .D(n283), .Z(N86) );
  GTECH_OAI2N2 U274 ( .A(n25), .B(n285), .C(R[2]), .D(n283), .Z(N85) );
  GTECH_OAI2N2 U275 ( .A(n26), .B(n285), .C(R[1]), .D(n283), .Z(N84) );
  GTECH_OAI2N2 U276 ( .A(n27), .B(n285), .C(R[0]), .D(n283), .Z(N83) );
  GTECH_NOT U277 ( .A(n286), .Z(N82) );
  GTECH_AND2 U278 ( .A(M[15]), .B(n283), .Z(N42) );
  GTECH_AND2 U279 ( .A(M[14]), .B(n283), .Z(N39) );
  GTECH_AND2 U280 ( .A(M[13]), .B(n283), .Z(N38) );
  GTECH_AND2 U281 ( .A(M[12]), .B(n283), .Z(N37) );
  GTECH_AND2 U282 ( .A(M[11]), .B(n283), .Z(N36) );
  GTECH_AND2 U283 ( .A(M[10]), .B(n283), .Z(N35) );
  GTECH_AND2 U284 ( .A(M[9]), .B(n283), .Z(N34) );
  GTECH_AND2 U285 ( .A(M[8]), .B(n283), .Z(N33) );
  GTECH_AND2 U286 ( .A(M[7]), .B(n283), .Z(N32) );
  GTECH_AND2 U287 ( .A(M[6]), .B(n283), .Z(N31) );
  GTECH_AND2 U288 ( .A(M[5]), .B(n283), .Z(N30) );
  GTECH_AND2 U289 ( .A(M[4]), .B(n283), .Z(N29) );
  GTECH_AND2 U290 ( .A(M[3]), .B(n283), .Z(N28) );
  GTECH_AND2 U291 ( .A(M[2]), .B(n283), .Z(N27) );
  GTECH_AND2 U292 ( .A(M[1]), .B(n283), .Z(N26) );
  GTECH_AND2 U293 ( .A(M[0]), .B(n283), .Z(N25) );
  GTECH_OAI21 U294 ( .A(n285), .B(n287), .C(n288), .Z(N19) );
  GTECH_OR_NOT U295 ( .A(n9), .B(n289), .Z(n287) );
  GTECH_NAND3 U296 ( .A(n290), .B(n291), .C(n285), .Z(N18) );
  GTECH_AOI21 U297 ( .A(n289), .B(n292), .C(n285), .Z(N17) );
  GTECH_OR_NOT U298 ( .A(n8), .B(n293), .Z(n292) );
  GTECH_AOI21 U299 ( .A(n293), .B(n294), .C(n285), .Z(N16) );
  GTECH_OR_NOT U300 ( .A(n7), .B(n295), .Z(n294) );
  GTECH_NOT U301 ( .A(n296), .Z(N152) );
  GTECH_AOI222 U302 ( .A(n297), .B(n298), .C(n299), .D(n300), .E(n301), .F(
        n302), .Z(n296) );
  GTECH_OR_NOT U303 ( .A(N155), .B(n291), .Z(N151) );
  GTECH_NOT U304 ( .A(n303), .Z(N150) );
  GTECH_AOI222 U305 ( .A(n304), .B(n297), .C(n299), .D(n305), .E(n306), .F(
        n301), .Z(n303) );
  GTECH_MUX2 U306 ( .A(n307), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND2 U307 ( .A(n308), .B(n309), .Z(n307) );
  GTECH_NOT U308 ( .A(n310), .Z(N149) );
  GTECH_AOI222 U309 ( .A(n311), .B(n297), .C(n299), .D(n312), .E(n313), .F(
        n301), .Z(n310) );
  GTECH_NOT U310 ( .A(n314), .Z(N148) );
  GTECH_AOI222 U311 ( .A(n315), .B(n297), .C(n299), .D(n316), .E(n317), .F(
        n301), .Z(n314) );
  GTECH_NOT U312 ( .A(n318), .Z(N147) );
  GTECH_AOI222 U313 ( .A(n319), .B(n297), .C(n299), .D(n320), .E(n321), .F(
        n301), .Z(n318) );
  GTECH_NOT U314 ( .A(n322), .Z(N146) );
  GTECH_AOI222 U315 ( .A(n323), .B(n297), .C(n299), .D(n324), .E(n325), .F(
        n301), .Z(n322) );
  GTECH_NOT U316 ( .A(n326), .Z(N145) );
  GTECH_AOI222 U317 ( .A(n327), .B(n297), .C(n299), .D(n328), .E(n329), .F(
        n301), .Z(n326) );
  GTECH_NOT U318 ( .A(n330), .Z(N144) );
  GTECH_AOI222 U319 ( .A(n331), .B(n297), .C(n299), .D(n332), .E(n333), .F(
        n301), .Z(n330) );
  GTECH_NOT U320 ( .A(n334), .Z(N143) );
  GTECH_AOI222 U321 ( .A(n335), .B(n297), .C(n299), .D(n336), .E(n337), .F(
        n301), .Z(n334) );
  GTECH_NOT U322 ( .A(n338), .Z(N142) );
  GTECH_AOI222 U323 ( .A(n339), .B(n297), .C(n299), .D(n340), .E(n341), .F(
        n301), .Z(n338) );
  GTECH_NOT U324 ( .A(n342), .Z(N141) );
  GTECH_AOI222 U325 ( .A(n343), .B(n297), .C(n299), .D(n344), .E(n345), .F(
        n301), .Z(n342) );
  GTECH_NOT U326 ( .A(n346), .Z(N140) );
  GTECH_AOI222 U327 ( .A(n347), .B(n297), .C(n299), .D(n348), .E(n349), .F(
        n301), .Z(n346) );
  GTECH_NOT U328 ( .A(n350), .Z(N14) );
  GTECH_OR_NOT U329 ( .A(n309), .B(n308), .Z(n350) );
  GTECH_NOT U330 ( .A(n351), .Z(N139) );
  GTECH_AOI222 U331 ( .A(n352), .B(n297), .C(n299), .D(n353), .E(n354), .F(
        n301), .Z(n351) );
  GTECH_NOT U332 ( .A(n355), .Z(N138) );
  GTECH_AOI222 U333 ( .A(n356), .B(n297), .C(n299), .D(n357), .E(n358), .F(
        n301), .Z(n355) );
  GTECH_NOT U334 ( .A(n359), .Z(N137) );
  GTECH_AOI222 U335 ( .A(n360), .B(n297), .C(n299), .D(n361), .E(n362), .F(
        n301), .Z(n359) );
  GTECH_NOT U336 ( .A(n363), .Z(N136) );
  GTECH_AOI222 U337 ( .A(n299), .B(n274), .C(n301), .D(n276), .E(n297), .F(
        n278), .Z(n363) );
  GTECH_NOT U338 ( .A(n364), .Z(n278) );
  GTECH_XOR2 U339 ( .A(n365), .B(n366), .Z(n364) );
  GTECH_NOT U340 ( .A(n367), .Z(n276) );
  GTECH_XOR2 U341 ( .A(n365), .B(n368), .Z(n367) );
  GTECH_XOR2 U342 ( .A(n274), .B(n256), .Z(n365) );
  GTECH_NOT U343 ( .A(n369), .Z(n299) );
  GTECH_OAI21 U344 ( .A(n12), .B(n369), .C(n370), .Z(N135) );
  GTECH_OAI21 U345 ( .A(n301), .B(n297), .C(n282), .Z(n370) );
  GTECH_OAI21 U346 ( .A(n12), .B(n371), .C(n372), .Z(n282) );
  GTECH_NOT U347 ( .A(n255), .Z(n371) );
  GTECH_NOT U348 ( .A(n373), .Z(n297) );
  GTECH_NAND3 U349 ( .A(n28), .B(n374), .C(N155), .Z(n373) );
  GTECH_NOT U350 ( .A(n375), .Z(n301) );
  GTECH_NAND3 U351 ( .A(n10), .B(n376), .C(N155), .Z(n375) );
  GTECH_NOT U352 ( .A(n28), .Z(n376) );
  GTECH_OR_NOT U353 ( .A(n377), .B(n378), .Z(n369) );
  GTECH_XOR2 U354 ( .A(n374), .B(n28), .Z(n378) );
  GTECH_AND2 U355 ( .A(N155), .B(n379), .Z(N134) );
  GTECH_NOT U356 ( .A(n13), .Z(n379) );
  GTECH_AND2 U357 ( .A(N155), .B(n380), .Z(N133) );
  GTECH_NOT U358 ( .A(n14), .Z(n380) );
  GTECH_AND2 U359 ( .A(N155), .B(n381), .Z(N132) );
  GTECH_NOT U360 ( .A(n15), .Z(n381) );
  GTECH_AND2 U361 ( .A(N155), .B(n382), .Z(N131) );
  GTECH_NOT U362 ( .A(n16), .Z(n382) );
  GTECH_AND2 U363 ( .A(N155), .B(n383), .Z(N130) );
  GTECH_NOT U364 ( .A(n17), .Z(n383) );
  GTECH_AND2 U365 ( .A(N155), .B(n384), .Z(N129) );
  GTECH_NOT U366 ( .A(n18), .Z(n384) );
  GTECH_AND2 U367 ( .A(N155), .B(n385), .Z(N128) );
  GTECH_NOT U368 ( .A(n19), .Z(n385) );
  GTECH_AND2 U369 ( .A(N155), .B(n386), .Z(N127) );
  GTECH_NOT U370 ( .A(n20), .Z(n386) );
  GTECH_AND2 U371 ( .A(N155), .B(n387), .Z(N126) );
  GTECH_NOT U372 ( .A(n21), .Z(n387) );
  GTECH_AND2 U373 ( .A(N155), .B(n388), .Z(N125) );
  GTECH_NOT U374 ( .A(n22), .Z(n388) );
  GTECH_AND2 U375 ( .A(N155), .B(n389), .Z(N124) );
  GTECH_NOT U376 ( .A(n23), .Z(n389) );
  GTECH_AND2 U377 ( .A(N155), .B(n390), .Z(N123) );
  GTECH_NOT U378 ( .A(n24), .Z(n390) );
  GTECH_AND2 U379 ( .A(N155), .B(n391), .Z(N122) );
  GTECH_NOT U380 ( .A(n25), .Z(n391) );
  GTECH_AND2 U381 ( .A(N155), .B(n392), .Z(N121) );
  GTECH_NOT U382 ( .A(n26), .Z(n392) );
  GTECH_AND2 U383 ( .A(N155), .B(n393), .Z(N120) );
  GTECH_NOT U384 ( .A(n27), .Z(n393) );
  GTECH_NOT U385 ( .A(n377), .Z(N155) );
  GTECH_NAND4 U386 ( .A(n8), .B(n7), .C(n9), .D(n394), .Z(n377) );
  GTECH_AND3 U387 ( .A(n291), .B(n309), .C(n6), .Z(n394) );
  GTECH_NOT U388 ( .A(n395), .Z(N116) );
  GTECH_AOI222 U389 ( .A(n273), .B(n300), .C(n302), .D(n275), .E(n298), .F(
        n277), .Z(n395) );
  GTECH_XOR2 U390 ( .A(n396), .B(n397), .Z(n298) );
  GTECH_OA21 U391 ( .A(n31), .B(n270), .C(n398), .Z(n397) );
  GTECH_OAI21 U392 ( .A(n399), .B(n305), .C(n400), .Z(n398) );
  GTECH_XOR2 U393 ( .A(n396), .B(n401), .Z(n302) );
  GTECH_OA21 U394 ( .A(n270), .B(n305), .C(n402), .Z(n401) );
  GTECH_OAI21 U395 ( .A(n31), .B(n399), .C(n403), .Z(n402) );
  GTECH_XOR2 U396 ( .A(A[16]), .B(n30), .Z(n396) );
  GTECH_NOT U397 ( .A(n30), .Z(n300) );
  GTECH_OR_NOT U398 ( .A(N41), .B(n285), .Z(N115) );
  GTECH_OR_NOT U399 ( .A(n283), .B(n291), .Z(N41) );
  GTECH_NOT U400 ( .A(n288), .Z(n283) );
  GTECH_OR_NOT U401 ( .A(Rst), .B(Ld), .Z(n288) );
  GTECH_NOT U402 ( .A(n404), .Z(N113) );
  GTECH_AOI222 U403 ( .A(n273), .B(n305), .C(n306), .D(n275), .E(n304), .F(
        n277), .Z(n404) );
  GTECH_XOR2 U404 ( .A(n405), .B(n406), .Z(n304) );
  GTECH_NOT U405 ( .A(n400), .Z(n406) );
  GTECH_OAI21 U406 ( .A(n32), .B(n269), .C(n407), .Z(n400) );
  GTECH_OAI21 U407 ( .A(n408), .B(n312), .C(n409), .Z(n407) );
  GTECH_XOR2 U408 ( .A(n405), .B(n410), .Z(n306) );
  GTECH_NOT U409 ( .A(n403), .Z(n410) );
  GTECH_OAI21 U410 ( .A(n269), .B(n312), .C(n411), .Z(n403) );
  GTECH_OAI21 U411 ( .A(n32), .B(n408), .C(n412), .Z(n411) );
  GTECH_XOR2 U412 ( .A(n399), .B(n31), .Z(n405) );
  GTECH_NOT U413 ( .A(n270), .Z(n399) );
  GTECH_NOT U414 ( .A(n31), .Z(n305) );
  GTECH_NOT U415 ( .A(n413), .Z(N112) );
  GTECH_AOI222 U416 ( .A(n273), .B(n312), .C(n313), .D(n275), .E(n311), .F(
        n277), .Z(n413) );
  GTECH_XOR2 U417 ( .A(n414), .B(n415), .Z(n311) );
  GTECH_NOT U418 ( .A(n409), .Z(n415) );
  GTECH_OAI21 U419 ( .A(n33), .B(n268), .C(n416), .Z(n409) );
  GTECH_OAI21 U420 ( .A(n417), .B(n316), .C(n418), .Z(n416) );
  GTECH_XOR2 U421 ( .A(n414), .B(n419), .Z(n313) );
  GTECH_NOT U422 ( .A(n412), .Z(n419) );
  GTECH_OAI21 U423 ( .A(n268), .B(n316), .C(n420), .Z(n412) );
  GTECH_OAI21 U424 ( .A(n33), .B(n417), .C(n421), .Z(n420) );
  GTECH_XOR2 U425 ( .A(n408), .B(n32), .Z(n414) );
  GTECH_NOT U426 ( .A(n269), .Z(n408) );
  GTECH_NOT U427 ( .A(n32), .Z(n312) );
  GTECH_NOT U428 ( .A(n422), .Z(N111) );
  GTECH_AOI222 U429 ( .A(n273), .B(n316), .C(n317), .D(n275), .E(n315), .F(
        n277), .Z(n422) );
  GTECH_XOR2 U430 ( .A(n423), .B(n424), .Z(n315) );
  GTECH_NOT U431 ( .A(n418), .Z(n424) );
  GTECH_OAI21 U432 ( .A(n34), .B(n267), .C(n425), .Z(n418) );
  GTECH_OAI21 U433 ( .A(n426), .B(n320), .C(n427), .Z(n425) );
  GTECH_XOR2 U434 ( .A(n423), .B(n428), .Z(n317) );
  GTECH_NOT U435 ( .A(n421), .Z(n428) );
  GTECH_OAI21 U436 ( .A(n267), .B(n320), .C(n429), .Z(n421) );
  GTECH_OAI21 U437 ( .A(n34), .B(n426), .C(n430), .Z(n429) );
  GTECH_XOR2 U438 ( .A(n417), .B(n33), .Z(n423) );
  GTECH_NOT U439 ( .A(n268), .Z(n417) );
  GTECH_NOT U440 ( .A(n33), .Z(n316) );
  GTECH_NOT U441 ( .A(n431), .Z(N110) );
  GTECH_AOI222 U442 ( .A(n273), .B(n320), .C(n321), .D(n275), .E(n319), .F(
        n277), .Z(n431) );
  GTECH_XOR2 U443 ( .A(n432), .B(n433), .Z(n319) );
  GTECH_NOT U444 ( .A(n427), .Z(n433) );
  GTECH_OAI21 U445 ( .A(n35), .B(n266), .C(n434), .Z(n427) );
  GTECH_OAI21 U446 ( .A(n435), .B(n324), .C(n436), .Z(n434) );
  GTECH_XOR2 U447 ( .A(n432), .B(n437), .Z(n321) );
  GTECH_NOT U448 ( .A(n430), .Z(n437) );
  GTECH_OAI21 U449 ( .A(n266), .B(n324), .C(n438), .Z(n430) );
  GTECH_OAI21 U450 ( .A(n35), .B(n435), .C(n439), .Z(n438) );
  GTECH_XOR2 U451 ( .A(n426), .B(n34), .Z(n432) );
  GTECH_NOT U452 ( .A(n267), .Z(n426) );
  GTECH_NOT U453 ( .A(n34), .Z(n320) );
  GTECH_NOT U454 ( .A(n440), .Z(N109) );
  GTECH_AOI222 U455 ( .A(n273), .B(n324), .C(n325), .D(n275), .E(n323), .F(
        n277), .Z(n440) );
  GTECH_XOR2 U456 ( .A(n441), .B(n442), .Z(n323) );
  GTECH_NOT U457 ( .A(n436), .Z(n442) );
  GTECH_OAI21 U458 ( .A(n36), .B(n265), .C(n443), .Z(n436) );
  GTECH_OAI21 U459 ( .A(n444), .B(n328), .C(n445), .Z(n443) );
  GTECH_XOR2 U460 ( .A(n441), .B(n446), .Z(n325) );
  GTECH_NOT U461 ( .A(n439), .Z(n446) );
  GTECH_OAI21 U462 ( .A(n265), .B(n328), .C(n447), .Z(n439) );
  GTECH_OAI21 U463 ( .A(n36), .B(n444), .C(n448), .Z(n447) );
  GTECH_XOR2 U464 ( .A(n435), .B(n35), .Z(n441) );
  GTECH_NOT U465 ( .A(n266), .Z(n435) );
  GTECH_NOT U466 ( .A(n35), .Z(n324) );
  GTECH_NOT U467 ( .A(n449), .Z(N108) );
  GTECH_AOI222 U468 ( .A(n273), .B(n328), .C(n329), .D(n275), .E(n327), .F(
        n277), .Z(n449) );
  GTECH_XOR2 U469 ( .A(n450), .B(n451), .Z(n327) );
  GTECH_NOT U470 ( .A(n445), .Z(n451) );
  GTECH_OAI21 U471 ( .A(n37), .B(n264), .C(n452), .Z(n445) );
  GTECH_OAI21 U472 ( .A(n453), .B(n332), .C(n454), .Z(n452) );
  GTECH_XOR2 U473 ( .A(n450), .B(n455), .Z(n329) );
  GTECH_NOT U474 ( .A(n448), .Z(n455) );
  GTECH_OAI21 U475 ( .A(n264), .B(n332), .C(n456), .Z(n448) );
  GTECH_OAI21 U476 ( .A(n37), .B(n453), .C(n457), .Z(n456) );
  GTECH_XOR2 U477 ( .A(n444), .B(n36), .Z(n450) );
  GTECH_NOT U478 ( .A(n265), .Z(n444) );
  GTECH_NOT U479 ( .A(n36), .Z(n328) );
  GTECH_NOT U480 ( .A(n458), .Z(N107) );
  GTECH_AOI222 U481 ( .A(n273), .B(n332), .C(n333), .D(n275), .E(n331), .F(
        n277), .Z(n458) );
  GTECH_XOR2 U482 ( .A(n459), .B(n460), .Z(n331) );
  GTECH_NOT U483 ( .A(n454), .Z(n460) );
  GTECH_OAI21 U484 ( .A(n38), .B(n263), .C(n461), .Z(n454) );
  GTECH_OAI21 U485 ( .A(n462), .B(n336), .C(n463), .Z(n461) );
  GTECH_XOR2 U486 ( .A(n459), .B(n464), .Z(n333) );
  GTECH_NOT U487 ( .A(n457), .Z(n464) );
  GTECH_OAI21 U488 ( .A(n263), .B(n336), .C(n465), .Z(n457) );
  GTECH_OAI21 U489 ( .A(n38), .B(n462), .C(n466), .Z(n465) );
  GTECH_XOR2 U490 ( .A(n453), .B(n37), .Z(n459) );
  GTECH_NOT U491 ( .A(n264), .Z(n453) );
  GTECH_NOT U492 ( .A(n37), .Z(n332) );
  GTECH_NOT U493 ( .A(n467), .Z(N106) );
  GTECH_AOI222 U494 ( .A(n273), .B(n336), .C(n337), .D(n275), .E(n335), .F(
        n277), .Z(n467) );
  GTECH_XOR2 U495 ( .A(n468), .B(n469), .Z(n335) );
  GTECH_NOT U496 ( .A(n463), .Z(n469) );
  GTECH_OAI21 U497 ( .A(n39), .B(n262), .C(n470), .Z(n463) );
  GTECH_OAI21 U498 ( .A(n471), .B(n340), .C(n472), .Z(n470) );
  GTECH_XOR2 U499 ( .A(n468), .B(n473), .Z(n337) );
  GTECH_NOT U500 ( .A(n466), .Z(n473) );
  GTECH_OAI21 U501 ( .A(n262), .B(n340), .C(n474), .Z(n466) );
  GTECH_OAI21 U502 ( .A(n39), .B(n471), .C(n475), .Z(n474) );
  GTECH_XOR2 U503 ( .A(n462), .B(n38), .Z(n468) );
  GTECH_NOT U504 ( .A(n263), .Z(n462) );
  GTECH_NOT U505 ( .A(n38), .Z(n336) );
  GTECH_NOT U506 ( .A(n476), .Z(N105) );
  GTECH_AOI222 U507 ( .A(n273), .B(n340), .C(n341), .D(n275), .E(n339), .F(
        n277), .Z(n476) );
  GTECH_XOR2 U508 ( .A(n477), .B(n478), .Z(n339) );
  GTECH_NOT U509 ( .A(n472), .Z(n478) );
  GTECH_OAI21 U510 ( .A(n40), .B(n261), .C(n479), .Z(n472) );
  GTECH_OAI21 U511 ( .A(n480), .B(n344), .C(n481), .Z(n479) );
  GTECH_XOR2 U512 ( .A(n477), .B(n482), .Z(n341) );
  GTECH_NOT U513 ( .A(n475), .Z(n482) );
  GTECH_OAI21 U514 ( .A(n261), .B(n344), .C(n483), .Z(n475) );
  GTECH_OAI21 U515 ( .A(n40), .B(n480), .C(n484), .Z(n483) );
  GTECH_XOR2 U516 ( .A(n471), .B(n39), .Z(n477) );
  GTECH_NOT U517 ( .A(n262), .Z(n471) );
  GTECH_NOT U518 ( .A(n39), .Z(n340) );
  GTECH_NOT U519 ( .A(n485), .Z(N104) );
  GTECH_AOI222 U520 ( .A(n273), .B(n344), .C(n345), .D(n275), .E(n343), .F(
        n277), .Z(n485) );
  GTECH_XOR2 U521 ( .A(n486), .B(n487), .Z(n343) );
  GTECH_NOT U522 ( .A(n481), .Z(n487) );
  GTECH_OAI21 U523 ( .A(n41), .B(n260), .C(n488), .Z(n481) );
  GTECH_OAI21 U524 ( .A(n489), .B(n348), .C(n490), .Z(n488) );
  GTECH_XOR2 U525 ( .A(n486), .B(n491), .Z(n345) );
  GTECH_NOT U526 ( .A(n484), .Z(n491) );
  GTECH_OAI21 U527 ( .A(n260), .B(n348), .C(n492), .Z(n484) );
  GTECH_OAI21 U528 ( .A(n41), .B(n489), .C(n493), .Z(n492) );
  GTECH_XOR2 U529 ( .A(n480), .B(n40), .Z(n486) );
  GTECH_NOT U530 ( .A(n261), .Z(n480) );
  GTECH_NOT U531 ( .A(n40), .Z(n344) );
  GTECH_NOT U532 ( .A(n494), .Z(N103) );
  GTECH_AOI222 U533 ( .A(n273), .B(n348), .C(n349), .D(n275), .E(n347), .F(
        n277), .Z(n494) );
  GTECH_XOR2 U534 ( .A(n495), .B(n496), .Z(n347) );
  GTECH_NOT U535 ( .A(n490), .Z(n496) );
  GTECH_OAI21 U536 ( .A(n42), .B(n259), .C(n497), .Z(n490) );
  GTECH_OAI21 U537 ( .A(n498), .B(n353), .C(n499), .Z(n497) );
  GTECH_XOR2 U538 ( .A(n495), .B(n500), .Z(n349) );
  GTECH_NOT U539 ( .A(n493), .Z(n500) );
  GTECH_OAI21 U540 ( .A(n259), .B(n353), .C(n501), .Z(n493) );
  GTECH_OAI21 U541 ( .A(n42), .B(n498), .C(n502), .Z(n501) );
  GTECH_XOR2 U542 ( .A(n489), .B(n41), .Z(n495) );
  GTECH_NOT U543 ( .A(n260), .Z(n489) );
  GTECH_NOT U544 ( .A(n41), .Z(n348) );
  GTECH_NOT U545 ( .A(n503), .Z(N102) );
  GTECH_AOI222 U546 ( .A(n273), .B(n353), .C(n354), .D(n275), .E(n352), .F(
        n277), .Z(n503) );
  GTECH_XOR2 U547 ( .A(n504), .B(n505), .Z(n352) );
  GTECH_NOT U548 ( .A(n499), .Z(n505) );
  GTECH_OAI21 U549 ( .A(n43), .B(n258), .C(n506), .Z(n499) );
  GTECH_OAI21 U550 ( .A(n507), .B(n357), .C(n508), .Z(n506) );
  GTECH_XOR2 U551 ( .A(n504), .B(n509), .Z(n354) );
  GTECH_NOT U552 ( .A(n502), .Z(n509) );
  GTECH_OAI21 U553 ( .A(n258), .B(n357), .C(n510), .Z(n502) );
  GTECH_OAI21 U554 ( .A(n43), .B(n507), .C(n511), .Z(n510) );
  GTECH_XOR2 U555 ( .A(n498), .B(n42), .Z(n504) );
  GTECH_NOT U556 ( .A(n259), .Z(n498) );
  GTECH_NOT U557 ( .A(n42), .Z(n353) );
  GTECH_NOT U558 ( .A(n512), .Z(N101) );
  GTECH_AOI222 U559 ( .A(n273), .B(n357), .C(n358), .D(n275), .E(n356), .F(
        n277), .Z(n512) );
  GTECH_XOR2 U560 ( .A(n513), .B(n514), .Z(n356) );
  GTECH_NOT U561 ( .A(n508), .Z(n514) );
  GTECH_OAI21 U562 ( .A(n29), .B(n257), .C(n515), .Z(n508) );
  GTECH_OAI21 U563 ( .A(n516), .B(n361), .C(n517), .Z(n515) );
  GTECH_XOR2 U564 ( .A(n513), .B(n518), .Z(n358) );
  GTECH_NOT U565 ( .A(n511), .Z(n518) );
  GTECH_OAI21 U566 ( .A(n257), .B(n361), .C(n519), .Z(n511) );
  GTECH_OAI21 U567 ( .A(n29), .B(n516), .C(n520), .Z(n519) );
  GTECH_XOR2 U568 ( .A(n507), .B(n43), .Z(n513) );
  GTECH_NOT U569 ( .A(n258), .Z(n507) );
  GTECH_NOT U570 ( .A(n43), .Z(n357) );
  GTECH_NOT U571 ( .A(n521), .Z(N100) );
  GTECH_AOI222 U572 ( .A(n360), .B(n277), .C(n273), .D(n361), .E(n362), .F(
        n275), .Z(n521) );
  GTECH_NOT U573 ( .A(n522), .Z(n275) );
  GTECH_OR_NOT U574 ( .A(n286), .B(n10), .Z(n522) );
  GTECH_XOR2 U575 ( .A(n523), .B(n524), .Z(n362) );
  GTECH_NOT U576 ( .A(n520), .Z(n524) );
  GTECH_OAI21 U577 ( .A(n256), .B(n274), .C(n525), .Z(n520) );
  GTECH_OAI21 U578 ( .A(n11), .B(n526), .C(n368), .Z(n525) );
  GTECH_NOT U579 ( .A(n372), .Z(n368) );
  GTECH_OR_NOT U580 ( .A(n255), .B(n12), .Z(n372) );
  GTECH_NOT U581 ( .A(n29), .Z(n361) );
  GTECH_NOT U582 ( .A(n527), .Z(n273) );
  GTECH_MUX2 U583 ( .A(n286), .B(n528), .S(n10), .Z(n527) );
  GTECH_OR_NOT U584 ( .A(n285), .B(n28), .Z(n528) );
  GTECH_OR_NOT U585 ( .A(n28), .B(n308), .Z(n286) );
  GTECH_NOT U586 ( .A(n284), .Z(n277) );
  GTECH_NAND3 U587 ( .A(n308), .B(n374), .C(n28), .Z(n284) );
  GTECH_NOT U588 ( .A(n10), .Z(n374) );
  GTECH_NOT U589 ( .A(n285), .Z(n308) );
  GTECH_NAND3 U590 ( .A(n290), .B(n291), .C(n529), .Z(n285) );
  GTECH_OR_NOT U591 ( .A(n289), .B(n9), .Z(n529) );
  GTECH_OR_NOT U592 ( .A(n293), .B(n8), .Z(n289) );
  GTECH_OR_NOT U593 ( .A(n295), .B(n7), .Z(n293) );
  GTECH_OR_NOT U594 ( .A(n309), .B(n6), .Z(n295) );
  GTECH_NOT U595 ( .A(n254), .Z(n309) );
  GTECH_NOT U596 ( .A(Rst), .Z(n291) );
  GTECH_NOT U597 ( .A(Ld), .Z(n290) );
  GTECH_XOR2 U598 ( .A(n523), .B(n530), .Z(n360) );
  GTECH_NOT U599 ( .A(n517), .Z(n530) );
  GTECH_OAI21 U600 ( .A(n256), .B(n11), .C(n531), .Z(n517) );
  GTECH_OAI21 U601 ( .A(n526), .B(n274), .C(n366), .Z(n531) );
  GTECH_NOT U602 ( .A(n532), .Z(n366) );
  GTECH_OR_NOT U603 ( .A(n255), .B(n280), .Z(n532) );
  GTECH_NOT U604 ( .A(n12), .Z(n280) );
  GTECH_NOT U605 ( .A(n11), .Z(n274) );
  GTECH_NOT U606 ( .A(n256), .Z(n526) );
  GTECH_XOR2 U607 ( .A(n516), .B(n29), .Z(n523) );
  GTECH_NOT U608 ( .A(n257), .Z(n516) );
endmodule

