
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140;

  GTECH_XOR2 U93 ( .A(n74), .B(n75), .Z(sum[9]) );
  GTECH_XNOR2 U94 ( .A(n76), .B(n77), .Z(sum[8]) );
  GTECH_XNOR2 U95 ( .A(n78), .B(n79), .Z(sum[7]) );
  GTECH_OA21 U96 ( .A(n80), .B(n81), .C(n82), .Z(n79) );
  GTECH_XOR2 U97 ( .A(n80), .B(n81), .Z(sum[6]) );
  GTECH_AOI22 U98 ( .A(b[5]), .B(a[5]), .C(n83), .D(n84), .Z(n80) );
  GTECH_XOR2 U99 ( .A(n84), .B(n83), .Z(sum[5]) );
  GTECH_OAI21 U100 ( .A(n85), .B(n86), .C(n87), .Z(n83) );
  GTECH_XOR2 U101 ( .A(n86), .B(n85), .Z(sum[4]) );
  GTECH_NOT U102 ( .A(n88), .Z(n86) );
  GTECH_XNOR2 U103 ( .A(n89), .B(n90), .Z(sum[3]) );
  GTECH_AOI21 U104 ( .A(n91), .B(n92), .C(n93), .Z(n90) );
  GTECH_XOR2 U105 ( .A(n91), .B(n92), .Z(sum[2]) );
  GTECH_AO22 U106 ( .A(b[1]), .B(a[1]), .C(n94), .D(n95), .Z(n91) );
  GTECH_XOR2 U107 ( .A(n95), .B(n94), .Z(sum[1]) );
  GTECH_AO22 U108 ( .A(n96), .B(cin), .C(a[0]), .D(b[0]), .Z(n94) );
  GTECH_XOR2 U109 ( .A(n97), .B(n98), .Z(sum[15]) );
  GTECH_OA21 U110 ( .A(n99), .B(n100), .C(n101), .Z(n98) );
  GTECH_XOR2 U111 ( .A(n99), .B(n100), .Z(sum[14]) );
  GTECH_AOI2N2 U112 ( .A(b[13]), .B(a[13]), .C(n102), .D(n103), .Z(n99) );
  GTECH_XOR2 U113 ( .A(n103), .B(n102), .Z(sum[13]) );
  GTECH_OA21 U114 ( .A(n104), .B(n105), .C(n106), .Z(n102) );
  GTECH_NOT U115 ( .A(cout), .Z(n104) );
  GTECH_XNOR2 U116 ( .A(n105), .B(cout), .Z(sum[12]) );
  GTECH_XNOR2 U117 ( .A(n107), .B(n108), .Z(sum[11]) );
  GTECH_AOI21 U118 ( .A(n109), .B(n110), .C(n111), .Z(n108) );
  GTECH_XOR2 U119 ( .A(n109), .B(n110), .Z(sum[10]) );
  GTECH_AO22 U120 ( .A(b[9]), .B(a[9]), .C(n75), .D(n74), .Z(n109) );
  GTECH_AO22 U121 ( .A(n112), .B(n76), .C(a[8]), .D(b[8]), .Z(n75) );
  GTECH_XNOR2 U122 ( .A(n113), .B(n96), .Z(sum[0]) );
  GTECH_OAI21 U123 ( .A(n77), .B(n114), .C(n115), .Z(cout) );
  GTECH_NOT U124 ( .A(n112), .Z(n77) );
  GTECH_OAI21 U125 ( .A(n85), .B(n116), .C(n117), .Z(n112) );
  GTECH_OA21 U126 ( .A(n118), .B(n113), .C(n119), .Z(n85) );
  GTECH_NOT U127 ( .A(cin), .Z(n113) );
  GTECH_NOR3 U128 ( .A(n114), .B(n118), .C(n116), .Z(Pm) );
  GTECH_NAND5 U129 ( .A(n89), .B(n95), .C(n96), .D(n120), .E(n92), .Z(n118) );
  GTECH_XOR2 U130 ( .A(a[0]), .B(b[0]), .Z(n96) );
  GTECH_OAI21 U131 ( .A(n121), .B(n114), .C(n115), .Z(Gm) );
  GTECH_AOI2N2 U132 ( .A(b[15]), .B(a[15]), .C(n122), .D(n97), .Z(n115) );
  GTECH_OA21 U133 ( .A(n123), .B(n100), .C(n101), .Z(n122) );
  GTECH_AOI2N2 U134 ( .A(b[13]), .B(a[13]), .C(n103), .D(n106), .Z(n123) );
  GTECH_OR4 U135 ( .A(n105), .B(n100), .C(n97), .D(n103), .Z(n114) );
  GTECH_XNOR2 U136 ( .A(a[13]), .B(b[13]), .Z(n103) );
  GTECH_XNOR2 U137 ( .A(a[15]), .B(b[15]), .Z(n97) );
  GTECH_OAI21 U138 ( .A(b[14]), .B(a[14]), .C(n101), .Z(n100) );
  GTECH_NAND2 U139 ( .A(b[14]), .B(a[14]), .Z(n101) );
  GTECH_OAI21 U140 ( .A(b[12]), .B(a[12]), .C(n106), .Z(n105) );
  GTECH_NAND2 U141 ( .A(a[12]), .B(b[12]), .Z(n106) );
  GTECH_OA21 U142 ( .A(n119), .B(n116), .C(n117), .Z(n121) );
  GTECH_AOI2N2 U143 ( .A(b[11]), .B(a[11]), .C(n124), .D(n125), .Z(n117) );
  GTECH_NOT U144 ( .A(n107), .Z(n125) );
  GTECH_AOI21 U145 ( .A(n126), .B(n110), .C(n111), .Z(n124) );
  GTECH_AO21 U146 ( .A(b[9]), .B(a[9]), .C(n127), .Z(n126) );
  GTECH_NOT U147 ( .A(n128), .Z(n127) );
  GTECH_NAND3 U148 ( .A(a[8]), .B(n74), .C(b[8]), .Z(n128) );
  GTECH_NAND4 U149 ( .A(n110), .B(n76), .C(n107), .D(n74), .Z(n116) );
  GTECH_XOR2 U150 ( .A(a[9]), .B(b[9]), .Z(n74) );
  GTECH_XOR2 U151 ( .A(a[11]), .B(b[11]), .Z(n107) );
  GTECH_XOR2 U152 ( .A(a[8]), .B(b[8]), .Z(n76) );
  GTECH_OA21 U153 ( .A(a[10]), .B(b[10]), .C(n129), .Z(n110) );
  GTECH_NOT U154 ( .A(n111), .Z(n129) );
  GTECH_AND2 U155 ( .A(a[10]), .B(b[10]), .Z(n111) );
  GTECH_AOI222 U156 ( .A(n120), .B(n130), .C(b[7]), .D(a[7]), .E(n78), .F(n131), .Z(n119) );
  GTECH_OAI21 U157 ( .A(n132), .B(n81), .C(n82), .Z(n131) );
  GTECH_NOT U158 ( .A(n133), .Z(n81) );
  GTECH_AOI2N2 U159 ( .A(b[5]), .B(a[5]), .C(n134), .D(n87), .Z(n132) );
  GTECH_OAI2N2 U160 ( .A(n135), .B(n136), .C(b[3]), .D(a[3]), .Z(n130) );
  GTECH_NOT U161 ( .A(n89), .Z(n136) );
  GTECH_XOR2 U162 ( .A(a[3]), .B(b[3]), .Z(n89) );
  GTECH_AOI21 U163 ( .A(n137), .B(n92), .C(n93), .Z(n135) );
  GTECH_OA21 U164 ( .A(a[2]), .B(b[2]), .C(n138), .Z(n92) );
  GTECH_NOT U165 ( .A(n93), .Z(n138) );
  GTECH_AND2 U166 ( .A(a[2]), .B(b[2]), .Z(n93) );
  GTECH_AO21 U167 ( .A(b[1]), .B(a[1]), .C(n139), .Z(n137) );
  GTECH_NOT U168 ( .A(n140), .Z(n139) );
  GTECH_NAND3 U169 ( .A(a[0]), .B(n95), .C(b[0]), .Z(n140) );
  GTECH_XOR2 U170 ( .A(a[1]), .B(b[1]), .Z(n95) );
  GTECH_AND4 U171 ( .A(n88), .B(n133), .C(n84), .D(n78), .Z(n120) );
  GTECH_XOR2 U172 ( .A(a[7]), .B(b[7]), .Z(n78) );
  GTECH_NOT U173 ( .A(n134), .Z(n84) );
  GTECH_XNOR2 U174 ( .A(a[5]), .B(b[5]), .Z(n134) );
  GTECH_OA21 U175 ( .A(a[6]), .B(b[6]), .C(n82), .Z(n133) );
  GTECH_NAND2 U176 ( .A(b[6]), .B(a[6]), .Z(n82) );
  GTECH_OA21 U177 ( .A(b[4]), .B(a[4]), .C(n87), .Z(n88) );
  GTECH_NAND2 U178 ( .A(a[4]), .B(b[4]), .Z(n87) );
endmodule

