
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391;

  GTECH_MUX2 U140 ( .A(n279), .B(n280), .S(n281), .Z(sum[9]) );
  GTECH_XOR2 U141 ( .A(n282), .B(n283), .Z(n280) );
  GTECH_XOR2 U142 ( .A(n283), .B(n284), .Z(n279) );
  GTECH_AOI21 U143 ( .A(a[9]), .B(b[9]), .C(n285), .Z(n283) );
  GTECH_NOT U144 ( .A(n286), .Z(n285) );
  GTECH_XNOR2 U145 ( .A(n287), .B(n288), .Z(sum[8]) );
  GTECH_MUX2 U146 ( .A(n289), .B(n290), .S(n291), .Z(sum[7]) );
  GTECH_XNOR2 U147 ( .A(n292), .B(n293), .Z(n290) );
  GTECH_AND2 U148 ( .A(n294), .B(n295), .Z(n293) );
  GTECH_AO21 U149 ( .A(n296), .B(n297), .C(n298), .Z(n294) );
  GTECH_XOR2 U150 ( .A(n292), .B(n299), .Z(n289) );
  GTECH_XOR2 U151 ( .A(a[7]), .B(b[7]), .Z(n292) );
  GTECH_OAI21 U152 ( .A(n300), .B(n295), .C(n301), .Z(sum[6]) );
  GTECH_MUX2 U153 ( .A(n302), .B(n303), .S(n296), .Z(n301) );
  GTECH_XNOR2 U154 ( .A(n297), .B(n300), .Z(n303) );
  GTECH_OR_NOT U155 ( .A(a[6]), .B(n300), .Z(n302) );
  GTECH_OA21 U156 ( .A(n304), .B(n291), .C(n298), .Z(n300) );
  GTECH_OA21 U157 ( .A(n305), .B(n306), .C(n307), .Z(n298) );
  GTECH_MUX2 U158 ( .A(n308), .B(n309), .S(n310), .Z(sum[5]) );
  GTECH_AND2 U159 ( .A(n307), .B(n311), .Z(n310) );
  GTECH_OAI21 U160 ( .A(a[4]), .B(n312), .C(n313), .Z(n309) );
  GTECH_AO21 U161 ( .A(n312), .B(a[4]), .C(b[4]), .Z(n313) );
  GTECH_OAI21 U162 ( .A(n314), .B(n291), .C(n306), .Z(n308) );
  GTECH_XNOR2 U163 ( .A(n312), .B(n315), .Z(sum[4]) );
  GTECH_MUX2 U164 ( .A(n316), .B(n317), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U165 ( .A(n318), .B(n319), .Z(n317) );
  GTECH_XNOR2 U166 ( .A(n318), .B(n320), .Z(n316) );
  GTECH_AND_NOT U167 ( .A(n321), .B(n322), .Z(n320) );
  GTECH_AO21 U168 ( .A(n323), .B(n324), .C(n325), .Z(n321) );
  GTECH_XOR2 U169 ( .A(a[3]), .B(b[3]), .Z(n318) );
  GTECH_MUX2 U170 ( .A(n326), .B(n327), .S(n328), .Z(sum[2]) );
  GTECH_MUX2 U171 ( .A(n329), .B(n330), .S(n325), .Z(n327) );
  GTECH_OA21 U172 ( .A(n331), .B(n332), .C(n333), .Z(n325) );
  GTECH_MUX2 U173 ( .A(n330), .B(n329), .S(n334), .Z(n326) );
  GTECH_AO21 U174 ( .A(n323), .B(n324), .C(n322), .Z(n329) );
  GTECH_XNOR2 U175 ( .A(n324), .B(b[2]), .Z(n330) );
  GTECH_MUX2 U176 ( .A(n335), .B(n336), .S(n337), .Z(sum[1]) );
  GTECH_AND2 U177 ( .A(n333), .B(n338), .Z(n337) );
  GTECH_AO21 U178 ( .A(n328), .B(n332), .C(n339), .Z(n336) );
  GTECH_OAI21 U179 ( .A(n339), .B(n328), .C(n332), .Z(n335) );
  GTECH_NOT U180 ( .A(cin), .Z(n328) );
  GTECH_MUX2 U181 ( .A(n340), .B(n341), .S(n342), .Z(sum[15]) );
  GTECH_XNOR2 U182 ( .A(n343), .B(n344), .Z(n341) );
  GTECH_XOR2 U183 ( .A(n343), .B(n345), .Z(n340) );
  GTECH_AND2 U184 ( .A(n346), .B(n347), .Z(n345) );
  GTECH_OAI21 U185 ( .A(b[14]), .B(a[14]), .C(n348), .Z(n346) );
  GTECH_XNOR2 U186 ( .A(a[15]), .B(b[15]), .Z(n343) );
  GTECH_OAI21 U187 ( .A(n349), .B(n347), .C(n350), .Z(sum[14]) );
  GTECH_MUX2 U188 ( .A(n351), .B(n352), .S(b[14]), .Z(n350) );
  GTECH_OR_NOT U189 ( .A(a[14]), .B(n349), .Z(n352) );
  GTECH_XOR2 U190 ( .A(a[14]), .B(n349), .Z(n351) );
  GTECH_AOI21 U191 ( .A(n353), .B(n342), .C(n348), .Z(n349) );
  GTECH_AO22 U192 ( .A(a[13]), .B(b[13]), .C(n354), .D(n355), .Z(n348) );
  GTECH_MUX2 U193 ( .A(n356), .B(n357), .S(n342), .Z(sum[13]) );
  GTECH_XOR2 U194 ( .A(n358), .B(n359), .Z(n357) );
  GTECH_XOR2 U195 ( .A(n359), .B(n355), .Z(n356) );
  GTECH_AOI21 U196 ( .A(a[13]), .B(b[13]), .C(n360), .Z(n359) );
  GTECH_NOT U197 ( .A(n354), .Z(n360) );
  GTECH_XNOR2 U198 ( .A(n342), .B(n361), .Z(sum[12]) );
  GTECH_MUX2 U199 ( .A(n362), .B(n363), .S(n288), .Z(sum[11]) );
  GTECH_XNOR2 U200 ( .A(n364), .B(n365), .Z(n363) );
  GTECH_AND2 U201 ( .A(n366), .B(n367), .Z(n365) );
  GTECH_OAI21 U202 ( .A(b[10]), .B(a[10]), .C(n368), .Z(n366) );
  GTECH_XOR2 U203 ( .A(n364), .B(n369), .Z(n362) );
  GTECH_XOR2 U204 ( .A(a[11]), .B(b[11]), .Z(n364) );
  GTECH_OAI21 U205 ( .A(n370), .B(n367), .C(n371), .Z(sum[10]) );
  GTECH_MUX2 U206 ( .A(n372), .B(n373), .S(b[10]), .Z(n371) );
  GTECH_OR_NOT U207 ( .A(a[10]), .B(n370), .Z(n373) );
  GTECH_XOR2 U208 ( .A(a[10]), .B(n370), .Z(n372) );
  GTECH_AOI21 U209 ( .A(n374), .B(n281), .C(n368), .Z(n370) );
  GTECH_AO22 U210 ( .A(a[9]), .B(b[9]), .C(n286), .D(n284), .Z(n368) );
  GTECH_XOR2 U211 ( .A(cin), .B(n375), .Z(sum[0]) );
  GTECH_NOT U212 ( .A(n376), .Z(cout) );
  GTECH_MUX2 U213 ( .A(n361), .B(n377), .S(n342), .Z(n376) );
  GTECH_MUX2 U214 ( .A(n287), .B(n378), .S(n281), .Z(n342) );
  GTECH_NOT U215 ( .A(n288), .Z(n281) );
  GTECH_MUX2 U216 ( .A(n379), .B(n315), .S(n291), .Z(n288) );
  GTECH_NOT U217 ( .A(n312), .Z(n291) );
  GTECH_MUX2 U218 ( .A(n375), .B(n380), .S(cin), .Z(n312) );
  GTECH_OA21 U219 ( .A(a[3]), .B(n319), .C(n381), .Z(n380) );
  GTECH_AO21 U220 ( .A(n319), .B(a[3]), .C(b[3]), .Z(n381) );
  GTECH_OR_NOT U221 ( .A(n322), .B(n382), .Z(n319) );
  GTECH_AO21 U222 ( .A(n324), .B(n323), .C(n383), .Z(n382) );
  GTECH_NOT U223 ( .A(n334), .Z(n383) );
  GTECH_OAI21 U224 ( .A(n331), .B(n339), .C(n333), .Z(n334) );
  GTECH_NAND2 U225 ( .A(a[1]), .B(b[1]), .Z(n333) );
  GTECH_NOT U226 ( .A(n384), .Z(n339) );
  GTECH_NOT U227 ( .A(n338), .Z(n331) );
  GTECH_OR2 U228 ( .A(a[1]), .B(b[1]), .Z(n338) );
  GTECH_NOT U229 ( .A(b[2]), .Z(n323) );
  GTECH_NOT U230 ( .A(a[2]), .Z(n324) );
  GTECH_AND2 U231 ( .A(a[2]), .B(b[2]), .Z(n322) );
  GTECH_AND2 U232 ( .A(n332), .B(n384), .Z(n375) );
  GTECH_OR2 U233 ( .A(b[0]), .B(a[0]), .Z(n384) );
  GTECH_NAND2 U234 ( .A(b[0]), .B(a[0]), .Z(n332) );
  GTECH_OR_NOT U235 ( .A(n314), .B(n306), .Z(n315) );
  GTECH_NAND2 U236 ( .A(b[4]), .B(a[4]), .Z(n306) );
  GTECH_AOI21 U237 ( .A(n299), .B(a[7]), .C(n385), .Z(n379) );
  GTECH_OA21 U238 ( .A(a[7]), .B(n299), .C(b[7]), .Z(n385) );
  GTECH_NAND2 U239 ( .A(n386), .B(n295), .Z(n299) );
  GTECH_OR_NOT U240 ( .A(n296), .B(a[6]), .Z(n295) );
  GTECH_AO21 U241 ( .A(n297), .B(n296), .C(n304), .Z(n386) );
  GTECH_OA21 U242 ( .A(n314), .B(n305), .C(n307), .Z(n304) );
  GTECH_NAND2 U243 ( .A(b[5]), .B(a[5]), .Z(n307) );
  GTECH_NOT U244 ( .A(n311), .Z(n305) );
  GTECH_OR2 U245 ( .A(b[5]), .B(a[5]), .Z(n311) );
  GTECH_AND_NOT U246 ( .A(n387), .B(a[4]), .Z(n314) );
  GTECH_NOT U247 ( .A(b[4]), .Z(n387) );
  GTECH_NOT U248 ( .A(b[6]), .Z(n296) );
  GTECH_NOT U249 ( .A(a[6]), .Z(n297) );
  GTECH_OA21 U250 ( .A(a[11]), .B(n369), .C(n388), .Z(n378) );
  GTECH_AO21 U251 ( .A(n369), .B(a[11]), .C(b[11]), .Z(n388) );
  GTECH_NAND2 U252 ( .A(n389), .B(n367), .Z(n369) );
  GTECH_NAND2 U253 ( .A(a[10]), .B(b[10]), .Z(n367) );
  GTECH_OAI21 U254 ( .A(a[10]), .B(b[10]), .C(n374), .Z(n389) );
  GTECH_AO22 U255 ( .A(a[9]), .B(b[9]), .C(n282), .D(n286), .Z(n374) );
  GTECH_OR2 U256 ( .A(a[9]), .B(b[9]), .Z(n286) );
  GTECH_AND_NOT U257 ( .A(n282), .B(n284), .Z(n287) );
  GTECH_AND2 U258 ( .A(b[8]), .B(a[8]), .Z(n284) );
  GTECH_OR2 U259 ( .A(a[8]), .B(b[8]), .Z(n282) );
  GTECH_AOI21 U260 ( .A(n344), .B(a[15]), .C(n390), .Z(n377) );
  GTECH_OA21 U261 ( .A(a[15]), .B(n344), .C(b[15]), .Z(n390) );
  GTECH_NAND2 U262 ( .A(n391), .B(n347), .Z(n344) );
  GTECH_NAND2 U263 ( .A(a[14]), .B(b[14]), .Z(n347) );
  GTECH_OAI21 U264 ( .A(a[14]), .B(b[14]), .C(n353), .Z(n391) );
  GTECH_AO22 U265 ( .A(n354), .B(n358), .C(a[13]), .D(b[13]), .Z(n353) );
  GTECH_OR2 U266 ( .A(a[13]), .B(b[13]), .Z(n354) );
  GTECH_OR_NOT U267 ( .A(n355), .B(n358), .Z(n361) );
  GTECH_OR2 U268 ( .A(b[12]), .B(a[12]), .Z(n358) );
  GTECH_AND2 U269 ( .A(a[12]), .B(b[12]), .Z(n355) );
endmodule

