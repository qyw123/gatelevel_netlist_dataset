
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160;

  GTECH_XOR2 U101 ( .A(n82), .B(n83), .Z(sum[9]) );
  GTECH_XOR2 U102 ( .A(n84), .B(n85), .Z(sum[8]) );
  GTECH_XNOR2 U103 ( .A(n86), .B(n87), .Z(sum[7]) );
  GTECH_OAI21 U104 ( .A(n88), .B(n89), .C(n90), .Z(n86) );
  GTECH_XOR2 U105 ( .A(n89), .B(n88), .Z(sum[6]) );
  GTECH_OA21 U106 ( .A(n91), .B(n92), .C(n93), .Z(n88) );
  GTECH_XOR2 U107 ( .A(n92), .B(n91), .Z(sum[5]) );
  GTECH_OA21 U108 ( .A(n94), .B(n95), .C(n96), .Z(n91) );
  GTECH_XOR2 U109 ( .A(n95), .B(n94), .Z(sum[4]) );
  GTECH_XNOR2 U110 ( .A(n97), .B(n98), .Z(sum[3]) );
  GTECH_OA21 U111 ( .A(n99), .B(n100), .C(n101), .Z(n98) );
  GTECH_XNOR2 U112 ( .A(n102), .B(n99), .Z(sum[2]) );
  GTECH_AOI21 U113 ( .A(n103), .B(n104), .C(n105), .Z(n99) );
  GTECH_XOR2 U114 ( .A(n104), .B(n103), .Z(sum[1]) );
  GTECH_AO22 U115 ( .A(a[0]), .B(b[0]), .C(n106), .D(cin), .Z(n103) );
  GTECH_XOR2 U116 ( .A(n107), .B(n108), .Z(sum[15]) );
  GTECH_OA21 U117 ( .A(n109), .B(n110), .C(n111), .Z(n108) );
  GTECH_XOR2 U118 ( .A(n110), .B(n109), .Z(sum[14]) );
  GTECH_OA21 U119 ( .A(n112), .B(n113), .C(n114), .Z(n109) );
  GTECH_XOR2 U120 ( .A(n113), .B(n112), .Z(sum[13]) );
  GTECH_OA21 U121 ( .A(n115), .B(n116), .C(n117), .Z(n112) );
  GTECH_XOR2 U122 ( .A(n115), .B(n116), .Z(sum[12]) );
  GTECH_NOT U123 ( .A(cout), .Z(n115) );
  GTECH_XNOR2 U124 ( .A(n118), .B(n119), .Z(sum[11]) );
  GTECH_OAI21 U125 ( .A(n120), .B(n121), .C(n122), .Z(n118) );
  GTECH_XOR2 U126 ( .A(n121), .B(n120), .Z(sum[10]) );
  GTECH_OA21 U127 ( .A(n83), .B(n82), .C(n123), .Z(n120) );
  GTECH_OA21 U128 ( .A(n85), .B(n84), .C(n124), .Z(n83) );
  GTECH_XOR2 U129 ( .A(cin), .B(n106), .Z(sum[0]) );
  GTECH_OAI21 U130 ( .A(n85), .B(n125), .C(n126), .Z(cout) );
  GTECH_OA21 U131 ( .A(n94), .B(n127), .C(n128), .Z(n85) );
  GTECH_OA21 U132 ( .A(n129), .B(n130), .C(n131), .Z(n94) );
  GTECH_OR3 U133 ( .A(n132), .B(n100), .C(n133), .Z(n130) );
  GTECH_NOT U134 ( .A(cin), .Z(n133) );
  GTECH_NAND3 U135 ( .A(n97), .B(n104), .C(n106), .Z(n129) );
  GTECH_NOR4 U136 ( .A(n127), .B(n132), .C(n125), .D(n134), .Z(Pm) );
  GTECH_NAND4 U137 ( .A(n102), .B(n106), .C(n97), .D(n104), .Z(n134) );
  GTECH_XOR2 U138 ( .A(a[0]), .B(b[0]), .Z(n106) );
  GTECH_OAI21 U139 ( .A(n135), .B(n125), .C(n126), .Z(Gm) );
  GTECH_AOI2N2 U140 ( .A(b[15]), .B(a[15]), .C(n136), .D(n107), .Z(n126) );
  GTECH_OA21 U141 ( .A(n137), .B(n110), .C(n111), .Z(n136) );
  GTECH_OA21 U142 ( .A(n113), .B(n117), .C(n114), .Z(n137) );
  GTECH_OR4 U143 ( .A(n116), .B(n110), .C(n113), .D(n107), .Z(n125) );
  GTECH_XNOR2 U144 ( .A(a[15]), .B(b[15]), .Z(n107) );
  GTECH_OAI21 U145 ( .A(b[13]), .B(a[13]), .C(n114), .Z(n113) );
  GTECH_NOT U146 ( .A(n138), .Z(n114) );
  GTECH_AND2 U147 ( .A(b[13]), .B(a[13]), .Z(n138) );
  GTECH_OAI21 U148 ( .A(b[14]), .B(a[14]), .C(n111), .Z(n110) );
  GTECH_NOT U149 ( .A(n139), .Z(n111) );
  GTECH_AND2 U150 ( .A(b[14]), .B(a[14]), .Z(n139) );
  GTECH_OAI21 U151 ( .A(b[12]), .B(a[12]), .C(n117), .Z(n116) );
  GTECH_NOT U152 ( .A(n140), .Z(n117) );
  GTECH_AND2 U153 ( .A(b[12]), .B(a[12]), .Z(n140) );
  GTECH_OA21 U154 ( .A(n131), .B(n127), .C(n128), .Z(n135) );
  GTECH_OA21 U155 ( .A(n141), .B(n119), .C(n142), .Z(n128) );
  GTECH_OA21 U156 ( .A(n143), .B(n121), .C(n122), .Z(n141) );
  GTECH_OA21 U157 ( .A(n124), .B(n82), .C(n123), .Z(n143) );
  GTECH_OR4 U158 ( .A(n84), .B(n119), .C(n121), .D(n82), .Z(n127) );
  GTECH_OAI21 U159 ( .A(b[9]), .B(a[9]), .C(n123), .Z(n82) );
  GTECH_NOT U160 ( .A(n144), .Z(n123) );
  GTECH_AND2 U161 ( .A(b[9]), .B(a[9]), .Z(n144) );
  GTECH_OAI21 U162 ( .A(b[10]), .B(a[10]), .C(n122), .Z(n121) );
  GTECH_NOT U163 ( .A(n145), .Z(n122) );
  GTECH_AND2 U164 ( .A(b[10]), .B(a[10]), .Z(n145) );
  GTECH_OAI21 U165 ( .A(b[11]), .B(a[11]), .C(n142), .Z(n119) );
  GTECH_NOT U166 ( .A(n146), .Z(n142) );
  GTECH_AND2 U167 ( .A(b[11]), .B(a[11]), .Z(n146) );
  GTECH_OAI21 U168 ( .A(b[8]), .B(a[8]), .C(n124), .Z(n84) );
  GTECH_NOT U169 ( .A(n147), .Z(n124) );
  GTECH_AND2 U170 ( .A(b[8]), .B(a[8]), .Z(n147) );
  GTECH_OA21 U171 ( .A(n148), .B(n132), .C(n149), .Z(n131) );
  GTECH_OA21 U172 ( .A(n150), .B(n87), .C(n151), .Z(n149) );
  GTECH_OA21 U173 ( .A(n152), .B(n89), .C(n90), .Z(n150) );
  GTECH_OA21 U174 ( .A(n92), .B(n96), .C(n93), .Z(n152) );
  GTECH_OR4 U175 ( .A(n95), .B(n87), .C(n89), .D(n92), .Z(n132) );
  GTECH_OAI21 U176 ( .A(b[5]), .B(a[5]), .C(n93), .Z(n92) );
  GTECH_NOT U177 ( .A(n153), .Z(n93) );
  GTECH_AND2 U178 ( .A(b[5]), .B(a[5]), .Z(n153) );
  GTECH_OAI21 U179 ( .A(b[6]), .B(a[6]), .C(n90), .Z(n89) );
  GTECH_NOT U180 ( .A(n154), .Z(n90) );
  GTECH_AND2 U181 ( .A(b[6]), .B(a[6]), .Z(n154) );
  GTECH_OAI21 U182 ( .A(b[7]), .B(a[7]), .C(n151), .Z(n87) );
  GTECH_NOT U183 ( .A(n155), .Z(n151) );
  GTECH_AND2 U184 ( .A(b[7]), .B(a[7]), .Z(n155) );
  GTECH_OAI21 U185 ( .A(b[4]), .B(a[4]), .C(n96), .Z(n95) );
  GTECH_NOT U186 ( .A(n156), .Z(n96) );
  GTECH_AND2 U187 ( .A(b[4]), .B(a[4]), .Z(n156) );
  GTECH_AOI21 U188 ( .A(b[3]), .B(a[3]), .C(n157), .Z(n148) );
  GTECH_OA21 U189 ( .A(n158), .B(n159), .C(n97), .Z(n157) );
  GTECH_XOR2 U190 ( .A(a[3]), .B(b[3]), .Z(n97) );
  GTECH_OA21 U191 ( .A(n160), .B(n105), .C(n102), .Z(n158) );
  GTECH_NOT U192 ( .A(n100), .Z(n102) );
  GTECH_OAI21 U193 ( .A(b[2]), .B(a[2]), .C(n101), .Z(n100) );
  GTECH_NOT U194 ( .A(n159), .Z(n101) );
  GTECH_AND2 U195 ( .A(b[2]), .B(a[2]), .Z(n159) );
  GTECH_AND2 U196 ( .A(b[1]), .B(a[1]), .Z(n105) );
  GTECH_AND3 U197 ( .A(a[0]), .B(n104), .C(b[0]), .Z(n160) );
  GTECH_XOR2 U198 ( .A(a[1]), .B(b[1]), .Z(n104) );
endmodule

