
module fraction_multiplier4 ( CLK, St, Mplier, Mcand, Product, Done );
  input [3:0] Mplier;
  input [3:0] Mcand;
  output [6:0] Product;
  input CLK, St;
  output Done;
  wire   A_3_, N40, N41, N42, N44, N46, N48, N50, N52, N54, N56, N57, N58, N63,
         n12, n13, n14, n15, n16, n17, n18, n19, n71, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136;
  wire   [2:0] State;

  GTECH_FD1 State_reg_0_ ( .D(N40), .CP(CLK), .Q(State[0]), .QN(n12) );
  GTECH_FD1 State_reg_2_ ( .D(N42), .CP(CLK), .Q(State[2]), .QN(n13) );
  GTECH_FD1 State_reg_1_ ( .D(N41), .CP(CLK), .Q(State[1]), .QN(n81) );
  GTECH_FJK1S B_reg_0_ ( .J(n71), .K(n71), .TI(N52), .TE(N57), .CP(CLK), .Q(
        Product[0]), .QN(n14) );
  GTECH_FJK1S A_reg_3_ ( .J(n71), .K(n71), .TI(N50), .TE(N63), .CP(CLK), .Q(
        A_3_), .QN(n15) );
  GTECH_FJK1S A_reg_0_ ( .J(n71), .K(n71), .TI(N44), .TE(N57), .CP(CLK), .Q(
        Product[4]), .QN(n80) );
  GTECH_FJK1S A_reg_1_ ( .J(n71), .K(n71), .TI(N46), .TE(N57), .CP(CLK), .Q(
        Product[5]), .QN(n79) );
  GTECH_FJK1S A_reg_2_ ( .J(n71), .K(n71), .TI(N48), .TE(N57), .CP(CLK), .Q(
        Product[6]), .QN(n16) );
  GTECH_FJK1S B_reg_3_ ( .J(n71), .K(n71), .TI(N58), .TE(N57), .CP(CLK), .Q(
        Product[3]), .QN(n17) );
  GTECH_FJK1S B_reg_2_ ( .J(n71), .K(n71), .TI(N56), .TE(N57), .CP(CLK), .Q(
        Product[2]), .QN(n18) );
  GTECH_FJK1S B_reg_1_ ( .J(n71), .K(n71), .TI(N54), .TE(N57), .CP(CLK), .Q(
        Product[1]), .QN(n19) );
  GTECH_ZERO U76 ( .Z(n71) );
  GTECH_AND_NOT U77 ( .A(N57), .B(n82), .Z(N63) );
  GTECH_NOT U78 ( .A(n83), .Z(N58) );
  GTECH_AOI222 U79 ( .A(Mplier[3]), .B(n84), .C(n85), .D(n86), .E(n87), .F(n88), .Z(n83) );
  GTECH_OAI21 U80 ( .A(Mcand[0]), .B(n89), .C(n90), .Z(n87) );
  GTECH_NOT U81 ( .A(n82), .Z(n90) );
  GTECH_AND_NOT U82 ( .A(n91), .B(n14), .Z(n85) );
  GTECH_AO21 U83 ( .A(n84), .B(St), .C(n91), .Z(N57) );
  GTECH_NOT U84 ( .A(n89), .Z(n91) );
  GTECH_OAI2N2 U85 ( .A(n17), .B(n89), .C(Mplier[2]), .D(n84), .Z(N56) );
  GTECH_OAI2N2 U86 ( .A(n18), .B(n89), .C(Mplier[1]), .D(n84), .Z(N54) );
  GTECH_OAI2N2 U87 ( .A(n19), .B(n89), .C(Mplier[0]), .D(n84), .Z(N52) );
  GTECH_OAI22 U88 ( .A(Mcand[3]), .B(n92), .C(n93), .D(n94), .Z(N50) );
  GTECH_OAI21 U89 ( .A(n95), .B(n96), .C(n97), .Z(N48) );
  GTECH_OAI21 U90 ( .A(n82), .B(n98), .C(n96), .Z(n97) );
  GTECH_AO22 U91 ( .A(n94), .B(n99), .C(n100), .D(Mcand[3]), .Z(n98) );
  GTECH_NOT U92 ( .A(n15), .Z(n96) );
  GTECH_AOI22 U93 ( .A(n94), .B(n100), .C(n99), .D(Mcand[3]), .Z(n95) );
  GTECH_AO22 U94 ( .A(n101), .B(n102), .C(n103), .D(n104), .Z(n99) );
  GTECH_OAI22 U95 ( .A(n101), .B(n105), .C(n103), .D(n106), .Z(n100) );
  GTECH_OA21 U96 ( .A(n107), .B(n108), .C(n109), .Z(n103) );
  GTECH_AO21 U97 ( .A(n108), .B(n107), .C(n110), .Z(n109) );
  GTECH_OA21 U98 ( .A(n111), .B(n108), .C(n112), .Z(n101) );
  GTECH_AO21 U99 ( .A(n108), .B(n111), .C(n16), .Z(n112) );
  GTECH_NOT U100 ( .A(Mcand[3]), .Z(n94) );
  GTECH_OAI21 U101 ( .A(n110), .B(n113), .C(n114), .Z(N46) );
  GTECH_OAI21 U102 ( .A(n82), .B(n115), .C(n110), .Z(n114) );
  GTECH_AO22 U103 ( .A(n108), .B(n116), .C(n117), .D(Mcand[2]), .Z(n115) );
  GTECH_AOI22 U104 ( .A(n108), .B(n117), .C(n116), .D(Mcand[2]), .Z(n113) );
  GTECH_OAI2N2 U105 ( .A(n118), .B(n106), .C(n111), .D(n102), .Z(n116) );
  GTECH_NOT U106 ( .A(n119), .Z(n111) );
  GTECH_OAI2N2 U107 ( .A(n107), .B(n106), .C(n119), .D(n102), .Z(n117) );
  GTECH_ADD_ABC U108 ( .A(Mcand[1]), .B(n120), .C(n121), .COUT(n119) );
  GTECH_AND_NOT U109 ( .A(Mcand[0]), .B(n80), .Z(n120) );
  GTECH_NOT U110 ( .A(n118), .Z(n107) );
  GTECH_ADD_ABC U111 ( .A(n122), .B(Mcand[1]), .C(n79), .COUT(n118) );
  GTECH_AND_NOT U112 ( .A(Mcand[0]), .B(n88), .Z(n122) );
  GTECH_NOT U113 ( .A(n80), .Z(n88) );
  GTECH_NOT U114 ( .A(Mcand[2]), .Z(n108) );
  GTECH_NOT U115 ( .A(n16), .Z(n110) );
  GTECH_OAI21 U116 ( .A(n121), .B(n123), .C(n124), .Z(N44) );
  GTECH_OAI21 U117 ( .A(n82), .B(n125), .C(n121), .Z(n124) );
  GTECH_AO22 U118 ( .A(n126), .B(Mcand[1]), .C(n127), .D(n128), .Z(n125) );
  GTECH_AND_NOT U119 ( .A(n14), .B(n89), .Z(n82) );
  GTECH_AND_NOT U120 ( .A(n92), .B(n129), .Z(n89) );
  GTECH_AOI22 U121 ( .A(Mcand[1]), .B(n128), .C(n127), .D(n126), .Z(n123) );
  GTECH_OAI2N2 U122 ( .A(n130), .B(n105), .C(n86), .D(n104), .Z(n126) );
  GTECH_NOT U123 ( .A(Mcand[1]), .Z(n127) );
  GTECH_OA21 U124 ( .A(n104), .B(n130), .C(n131), .Z(n128) );
  GTECH_OAI21 U125 ( .A(n86), .B(n106), .C(n105), .Z(n131) );
  GTECH_NOT U126 ( .A(n102), .Z(n105) );
  GTECH_AND_NOT U127 ( .A(n129), .B(n14), .Z(n102) );
  GTECH_AND2 U128 ( .A(Mcand[0]), .B(n80), .Z(n86) );
  GTECH_OR_NOT U129 ( .A(n80), .B(Mcand[0]), .Z(n130) );
  GTECH_NOT U130 ( .A(n106), .Z(n104) );
  GTECH_OR2 U131 ( .A(n14), .B(n92), .Z(n106) );
  GTECH_NOT U132 ( .A(n79), .Z(n121) );
  GTECH_NAND2 U133 ( .A(n132), .B(n92), .Z(N42) );
  GTECH_OR3 U134 ( .A(n81), .B(n12), .C(n93), .Z(n132) );
  GTECH_OA21 U135 ( .A(n12), .B(n81), .C(n129), .Z(N41) );
  GTECH_AO21 U136 ( .A(n84), .B(St), .C(n133), .Z(N40) );
  GTECH_OAI21 U137 ( .A(n134), .B(n93), .C(n92), .Z(n133) );
  GTECH_OR_NOT U138 ( .A(n13), .B(n135), .Z(n92) );
  GTECH_NOT U139 ( .A(n129), .Z(n93) );
  GTECH_AND_NOT U140 ( .A(n13), .B(n135), .Z(n129) );
  GTECH_AND_NOT U141 ( .A(n135), .B(n136), .Z(n84) );
  GTECH_AND2 U142 ( .A(n81), .B(n12), .Z(n135) );
  GTECH_AND3 U143 ( .A(n134), .B(n136), .C(n81), .Z(Done) );
  GTECH_NOT U144 ( .A(n13), .Z(n136) );
  GTECH_NOT U145 ( .A(n12), .Z(n134) );
endmodule

