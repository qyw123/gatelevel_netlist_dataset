
module clock_12h ( clk, reset, ena, pm, hh, mm, ss );
  output [7:0] hh;
  output [7:0] mm;
  output [7:0] ss;
  input clk, reset, ena;
  output pm;
  wire   N22, N23, N24, N25, N26, N39, N40, N41, N42, N43, N55, N56, N57, N58,
         N59, N71, N72, N73, N74, N75, N88, N89, N90, N91, N92, N110, N112,
         N114, N115, N116, N121, N122, n4, n5, n6, n7, n8, n9, n10, n11, n85,
         n110, n111, n112, n113, n114, n115, n116, n117, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215;

  GTECH_FJK1S ss_ones_reg_0_ ( .J(n85), .K(n85), .TI(N22), .TE(N25), .CP(clk), 
        .Q(ss[0]) );
  GTECH_FJK1S ss_ones_reg_3_ ( .J(n85), .K(n85), .TI(N26), .TE(N25), .CP(clk), 
        .Q(ss[3]) );
  GTECH_FJK1S ss_ones_reg_1_ ( .J(n85), .K(n85), .TI(N23), .TE(N25), .CP(clk), 
        .Q(ss[1]) );
  GTECH_FJK1S ss_ones_reg_2_ ( .J(n85), .K(n85), .TI(N24), .TE(N25), .CP(clk), 
        .Q(ss[2]) );
  GTECH_FJK1S ss_tens_reg_0_ ( .J(n85), .K(n85), .TI(N39), .TE(N42), .CP(clk), 
        .Q(ss[4]) );
  GTECH_FJK1S ss_tens_reg_1_ ( .J(n85), .K(n85), .TI(N40), .TE(N42), .CP(clk), 
        .Q(ss[5]) );
  GTECH_FJK1S ss_tens_reg_2_ ( .J(n85), .K(n85), .TI(N41), .TE(N42), .CP(clk), 
        .Q(ss[6]) );
  GTECH_FJK1S ss_tens_reg_3_ ( .J(n85), .K(n85), .TI(N43), .TE(N42), .CP(clk), 
        .Q(ss[7]) );
  GTECH_FJK1S mm_ones_reg_0_ ( .J(n85), .K(n85), .TI(N55), .TE(N58), .CP(clk), 
        .Q(mm[0]), .QN(n4) );
  GTECH_FJK1S mm_ones_reg_3_ ( .J(n85), .K(n85), .TI(N59), .TE(N58), .CP(clk), 
        .Q(mm[3]), .QN(n115) );
  GTECH_FJK1S mm_ones_reg_1_ ( .J(n85), .K(n85), .TI(N56), .TE(N58), .CP(clk), 
        .Q(mm[1]), .QN(n117) );
  GTECH_FJK1S mm_ones_reg_2_ ( .J(n85), .K(n85), .TI(N57), .TE(N58), .CP(clk), 
        .Q(mm[2]), .QN(n116) );
  GTECH_FJK1S mm_tens_reg_0_ ( .J(n85), .K(n85), .TI(N71), .TE(N74), .CP(clk), 
        .Q(mm[4]), .QN(n114) );
  GTECH_FJK1S mm_tens_reg_1_ ( .J(n85), .K(n85), .TI(N72), .TE(N74), .CP(clk), 
        .Q(mm[5]), .QN(n113) );
  GTECH_FJK1S mm_tens_reg_2_ ( .J(n85), .K(n85), .TI(N73), .TE(N74), .CP(clk), 
        .Q(mm[6]), .QN(n112) );
  GTECH_FJK1S mm_tens_reg_3_ ( .J(n85), .K(n85), .TI(N75), .TE(N74), .CP(clk), 
        .Q(mm[7]), .QN(n5) );
  GTECH_FJK1S hh_tens_reg_0_ ( .J(n85), .K(n85), .TI(N110), .TE(N115), .CP(clk), .Q(hh[4]), .QN(n124) );
  GTECH_FJK1S hh_tens_reg_1_ ( .J(n85), .K(n85), .TI(N112), .TE(N115), .CP(clk), .Q(hh[5]), .QN(n6) );
  GTECH_FJK1S hh_tens_reg_2_ ( .J(n85), .K(n85), .TI(N114), .TE(N115), .CP(clk), .Q(hh[6]), .QN(n7) );
  GTECH_FJK1S hh_tens_reg_3_ ( .J(n85), .K(n85), .TI(N116), .TE(N115), .CP(clk), .Q(hh[7]), .QN(n8) );
  GTECH_FJK1S hh_ones_reg_0_ ( .J(n85), .K(n85), .TI(N88), .TE(N91), .CP(clk), 
        .Q(hh[0]), .QN(n9) );
  GTECH_FJK1S hh_ones_reg_1_ ( .J(n85), .K(n85), .TI(N89), .TE(N91), .CP(clk), 
        .Q(hh[1]), .QN(n111) );
  GTECH_FJK1S hh_ones_reg_2_ ( .J(n85), .K(n85), .TI(N90), .TE(N91), .CP(clk), 
        .Q(hh[2]), .QN(n10) );
  GTECH_FJK1S hh_ones_reg_3_ ( .J(n85), .K(n85), .TI(N92), .TE(N91), .CP(clk), 
        .Q(hh[3]), .QN(n110) );
  GTECH_FJK1S pm_temp_reg ( .J(n85), .K(n85), .TI(N122), .TE(N121), .CP(clk), 
        .Q(pm), .QN(n11) );
  GTECH_ZERO U133 ( .Z(n85) );
  GTECH_AND2 U134 ( .A(n125), .B(n126), .Z(N92) );
  GTECH_XOR2 U135 ( .A(n127), .B(n110), .Z(n125) );
  GTECH_OR2 U136 ( .A(n10), .B(n128), .Z(n127) );
  GTECH_NAND2 U137 ( .A(n129), .B(n130), .Z(N91) );
  GTECH_AND2 U138 ( .A(n131), .B(n126), .Z(N90) );
  GTECH_NOT U139 ( .A(n132), .Z(n126) );
  GTECH_XOR2 U140 ( .A(n128), .B(n10), .Z(n131) );
  GTECH_NAND2 U141 ( .A(n133), .B(n134), .Z(n128) );
  GTECH_OAI21 U142 ( .A(n135), .B(n132), .C(n129), .Z(N89) );
  GTECH_XOR2 U143 ( .A(n134), .B(n9), .Z(n135) );
  GTECH_OAI22 U144 ( .A(n130), .B(n136), .C(n133), .D(n132), .Z(N88) );
  GTECH_OR3 U145 ( .A(n137), .B(n138), .C(n130), .Z(n132) );
  GTECH_OAI22 U146 ( .A(n112), .B(n139), .C(n5), .D(n140), .Z(N75) );
  GTECH_OA21 U147 ( .A(n141), .B(n142), .C(n143), .Z(n140) );
  GTECH_OR_NOT U148 ( .A(n144), .B(n5), .Z(n139) );
  GTECH_OAI21 U149 ( .A(n112), .B(n143), .C(n145), .Z(N73) );
  GTECH_OR3 U150 ( .A(n113), .B(n144), .C(n141), .Z(n145) );
  GTECH_NOT U151 ( .A(n146), .Z(n143) );
  GTECH_OAI21 U152 ( .A(n147), .B(n142), .C(n148), .Z(n146) );
  GTECH_OAI22 U153 ( .A(n147), .B(n144), .C(n113), .D(n148), .Z(N72) );
  GTECH_NAND2 U154 ( .A(n149), .B(n150), .Z(n144) );
  GTECH_NOT U155 ( .A(n113), .Z(n147) );
  GTECH_NOT U156 ( .A(n148), .Z(N71) );
  GTECH_NAND2 U157 ( .A(n114), .B(n149), .Z(n148) );
  GTECH_NOT U158 ( .A(n142), .Z(n149) );
  GTECH_OR3 U159 ( .A(reset), .B(n151), .C(n152), .Z(n142) );
  GTECH_OAI22 U160 ( .A(n115), .B(n153), .C(n154), .D(n155), .Z(N59) );
  GTECH_OAI21 U161 ( .A(n116), .B(n115), .C(n156), .Z(n155) );
  GTECH_OAI21 U162 ( .A(n116), .B(n157), .C(n115), .Z(n156) );
  GTECH_OAI22 U163 ( .A(n157), .B(n158), .C(n116), .D(n153), .Z(N57) );
  GTECH_NAND2 U164 ( .A(n159), .B(n157), .Z(n153) );
  GTECH_OR_NOT U165 ( .A(n154), .B(n116), .Z(n158) );
  GTECH_NAND2 U166 ( .A(n160), .B(n161), .Z(n157) );
  GTECH_OAI21 U167 ( .A(n117), .B(n162), .C(n163), .Z(N56) );
  GTECH_OR3 U168 ( .A(n4), .B(n154), .C(n160), .Z(n163) );
  GTECH_NOT U169 ( .A(n117), .Z(n160) );
  GTECH_NOT U170 ( .A(n162), .Z(N55) );
  GTECH_NAND2 U171 ( .A(n4), .B(n159), .Z(n162) );
  GTECH_NOT U172 ( .A(n154), .Z(n159) );
  GTECH_NAND2 U173 ( .A(n164), .B(n165), .Z(n154) );
  GTECH_NOT U174 ( .A(N74), .Z(n165) );
  GTECH_NAND2 U175 ( .A(n129), .B(n152), .Z(N74) );
  GTECH_OAI21 U176 ( .A(n166), .B(n167), .C(n168), .Z(N43) );
  GTECH_OR3 U177 ( .A(n169), .B(n170), .C(ss[7]), .Z(n168) );
  GTECH_OA21 U178 ( .A(ss[6]), .B(n171), .C(n172), .Z(n166) );
  GTECH_OAI21 U179 ( .A(n172), .B(n169), .C(n173), .Z(N41) );
  GTECH_OR3 U180 ( .A(n170), .B(n174), .C(ss[6]), .Z(n173) );
  GTECH_NOT U181 ( .A(ss[6]), .Z(n169) );
  GTECH_NOT U182 ( .A(n175), .Z(n172) );
  GTECH_OAI21 U183 ( .A(ss[5]), .B(n171), .C(n176), .Z(n175) );
  GTECH_OAI22 U184 ( .A(n174), .B(n176), .C(ss[5]), .D(n170), .Z(N40) );
  GTECH_NAND2 U185 ( .A(n177), .B(ss[4]), .Z(n170) );
  GTECH_NOT U186 ( .A(n176), .Z(N39) );
  GTECH_NAND2 U187 ( .A(n177), .B(n178), .Z(n176) );
  GTECH_NOT U188 ( .A(ss[4]), .Z(n178) );
  GTECH_NOT U189 ( .A(n171), .Z(n177) );
  GTECH_NAND2 U190 ( .A(n179), .B(n180), .Z(n171) );
  GTECH_NOT U191 ( .A(N58), .Z(n180) );
  GTECH_NAND2 U192 ( .A(n129), .B(n181), .Z(N58) );
  GTECH_OAI2N2 U193 ( .A(n182), .B(n183), .C(ss[3]), .D(n184), .Z(N26) );
  GTECH_OAI21 U194 ( .A(n185), .B(ss[2]), .C(n186), .Z(n184) );
  GTECH_OR_NOT U195 ( .A(ss[3]), .B(ss[2]), .Z(n183) );
  GTECH_NAND2 U196 ( .A(n129), .B(n187), .Z(N25) );
  GTECH_NOT U197 ( .A(ena), .Z(n187) );
  GTECH_OAI22 U198 ( .A(n186), .B(n188), .C(ss[2]), .D(n182), .Z(N24) );
  GTECH_OR3 U199 ( .A(n189), .B(n185), .C(n190), .Z(n182) );
  GTECH_NOT U200 ( .A(n191), .Z(n186) );
  GTECH_OAI21 U201 ( .A(ss[1]), .B(n185), .C(n192), .Z(n191) );
  GTECH_OAI21 U202 ( .A(n190), .B(n192), .C(n193), .Z(N23) );
  GTECH_OR3 U203 ( .A(n189), .B(n185), .C(ss[1]), .Z(n193) );
  GTECH_NOT U204 ( .A(n192), .Z(N22) );
  GTECH_NAND2 U205 ( .A(n194), .B(n189), .Z(n192) );
  GTECH_NOT U206 ( .A(ss[0]), .Z(n189) );
  GTECH_NOT U207 ( .A(n185), .Z(n194) );
  GTECH_NAND2 U208 ( .A(ena), .B(n195), .Z(n185) );
  GTECH_NOT U209 ( .A(N42), .Z(n195) );
  GTECH_NAND2 U210 ( .A(n129), .B(n196), .Z(N42) );
  GTECH_AND2 U211 ( .A(n197), .B(n11), .Z(N122) );
  GTECH_NOT U212 ( .A(n198), .Z(n197) );
  GTECH_NAND2 U213 ( .A(n129), .B(n198), .Z(N121) );
  GTECH_NAND5 U214 ( .A(n199), .B(n8), .C(n7), .D(n6), .E(n200), .Z(n198) );
  GTECH_AND5 U215 ( .A(n201), .B(n133), .C(n10), .D(n110), .E(n111), .Z(n200)
         );
  GTECH_AND2 U216 ( .A(n202), .B(n203), .Z(N116) );
  GTECH_XOR2 U217 ( .A(n204), .B(n8), .Z(n202) );
  GTECH_OR2 U218 ( .A(n7), .B(n205), .Z(n204) );
  GTECH_OR3 U219 ( .A(reset), .B(n137), .C(n138), .Z(N115) );
  GTECH_NOT U220 ( .A(n136), .Z(n138) );
  GTECH_NAND5 U221 ( .A(n9), .B(n8), .C(n7), .D(n6), .E(n206), .Z(n136) );
  GTECH_AND5 U222 ( .A(n134), .B(n201), .C(n151), .D(n110), .E(n10), .Z(n206)
         );
  GTECH_NOT U223 ( .A(n111), .Z(n134) );
  GTECH_AND2 U224 ( .A(n207), .B(n203), .Z(N114) );
  GTECH_XOR2 U225 ( .A(n205), .B(n7), .Z(n207) );
  GTECH_NAND2 U226 ( .A(n208), .B(n201), .Z(n205) );
  GTECH_NOT U227 ( .A(n6), .Z(n208) );
  GTECH_AND2 U228 ( .A(n203), .B(n209), .Z(N112) );
  GTECH_XOR2 U229 ( .A(n6), .B(n124), .Z(n209) );
  GTECH_NOT U230 ( .A(n210), .Z(n203) );
  GTECH_OAI21 U231 ( .A(n210), .B(n201), .C(n129), .Z(N110) );
  GTECH_NOT U232 ( .A(n124), .Z(n201) );
  GTECH_NAND2 U233 ( .A(n137), .B(n199), .Z(n210) );
  GTECH_NOT U234 ( .A(n130), .Z(n199) );
  GTECH_NAND2 U235 ( .A(n151), .B(n129), .Z(n130) );
  GTECH_NOT U236 ( .A(reset), .Z(n129) );
  GTECH_NOT U237 ( .A(n211), .Z(n137) );
  GTECH_NAND5 U238 ( .A(n212), .B(n133), .C(n151), .D(n111), .E(n10), .Z(n211)
         );
  GTECH_NOT U239 ( .A(n213), .Z(n151) );
  GTECH_NAND5 U240 ( .A(n141), .B(n150), .C(n214), .D(n5), .E(n113), .Z(n213)
         );
  GTECH_NOT U241 ( .A(n152), .Z(n214) );
  GTECH_NAND5 U242 ( .A(n215), .B(n161), .C(n164), .D(n117), .E(n116), .Z(n152) );
  GTECH_NOT U243 ( .A(n181), .Z(n164) );
  GTECH_NAND5 U244 ( .A(n174), .B(n167), .C(n179), .D(ss[6]), .E(ss[4]), .Z(
        n181) );
  GTECH_NOT U245 ( .A(n196), .Z(n179) );
  GTECH_NAND5 U246 ( .A(n190), .B(n188), .C(ena), .D(ss[3]), .E(ss[0]), .Z(
        n196) );
  GTECH_NOT U247 ( .A(ss[2]), .Z(n188) );
  GTECH_NOT U248 ( .A(ss[1]), .Z(n190) );
  GTECH_NOT U249 ( .A(ss[7]), .Z(n167) );
  GTECH_NOT U250 ( .A(ss[5]), .Z(n174) );
  GTECH_NOT U251 ( .A(n4), .Z(n161) );
  GTECH_NOT U252 ( .A(n115), .Z(n215) );
  GTECH_NOT U253 ( .A(n114), .Z(n150) );
  GTECH_NOT U254 ( .A(n112), .Z(n141) );
  GTECH_NOT U255 ( .A(n9), .Z(n133) );
  GTECH_NOT U256 ( .A(n110), .Z(n212) );
endmodule

