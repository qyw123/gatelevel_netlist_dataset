
module CRC32 ( crcIn, data, crcOut );
  input [31:0] crcIn;
  input [7:0] data;
  output [31:0] crcOut;
  wire   n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54;

  GTECH_XOR2 U60 ( .A(crcIn[17]), .B(n28), .Z(crcOut[9]) );
  GTECH_XOR3 U61 ( .A(crcIn[16]), .B(n29), .C(n30), .Z(crcOut[8]) );
  GTECH_XOR3 U62 ( .A(crcIn[15]), .B(n31), .C(n32), .Z(crcOut[7]) );
  GTECH_XOR2 U63 ( .A(crcIn[14]), .B(n33), .Z(crcOut[6]) );
  GTECH_XOR3 U64 ( .A(crcIn[13]), .B(n34), .C(crcOut[31]), .Z(crcOut[5]) );
  GTECH_XOR3 U65 ( .A(crcIn[12]), .B(n31), .C(n35), .Z(crcOut[4]) );
  GTECH_NOT U66 ( .A(n36), .Z(crcOut[3]) );
  GTECH_XOR3 U67 ( .A(crcIn[11]), .B(n37), .C(n38), .Z(n36) );
  GTECH_XOR3 U68 ( .A(crcIn[10]), .B(n39), .C(n40), .Z(crcOut[2]) );
  GTECH_XOR2 U69 ( .A(n32), .B(crcOut[30]), .Z(crcOut[29]) );
  GTECH_XOR2 U70 ( .A(n31), .B(n33), .Z(crcOut[28]) );
  GTECH_XOR2 U71 ( .A(n41), .B(n42), .Z(n31) );
  GTECH_XOR3 U72 ( .A(n33), .B(n43), .C(crcOut[31]), .Z(crcOut[27]) );
  GTECH_XOR2 U73 ( .A(n44), .B(n28), .Z(crcOut[31]) );
  GTECH_XOR3 U74 ( .A(n39), .B(n35), .C(crcOut[30]), .Z(crcOut[26]) );
  GTECH_XOR2 U75 ( .A(n40), .B(n45), .Z(crcOut[30]) );
  GTECH_XOR2 U76 ( .A(n40), .B(n46), .Z(crcOut[25]) );
  GTECH_XOR2 U77 ( .A(n41), .B(n47), .Z(crcOut[24]) );
  GTECH_XOR2 U78 ( .A(crcIn[31]), .B(n48), .Z(crcOut[23]) );
  GTECH_XOR2 U79 ( .A(crcIn[30]), .B(n46), .Z(crcOut[22]) );
  GTECH_XOR3 U80 ( .A(n42), .B(n32), .C(n35), .Z(n46) );
  GTECH_XOR2 U81 ( .A(crcIn[29]), .B(n47), .Z(crcOut[21]) );
  GTECH_XOR3 U82 ( .A(n28), .B(n33), .C(n37), .Z(n47) );
  GTECH_XOR2 U83 ( .A(crcIn[28]), .B(n48), .Z(crcOut[20]) );
  GTECH_XOR2 U84 ( .A(n34), .B(n45), .Z(n48) );
  GTECH_XOR2 U85 ( .A(n43), .B(n39), .Z(n34) );
  GTECH_XOR3 U86 ( .A(crcIn[9]), .B(n41), .C(n43), .Z(crcOut[1]) );
  GTECH_XOR4 U87 ( .A(n35), .B(n38), .C(crcIn[27]), .D(n29), .Z(crcOut[19]) );
  GTECH_NOT U88 ( .A(n45), .Z(n29) );
  GTECH_XOR2 U89 ( .A(n49), .B(n50), .Z(n45) );
  GTECH_NOT U90 ( .A(n28), .Z(n50) );
  GTECH_XOR2 U91 ( .A(n32), .B(n30), .Z(n38) );
  GTECH_NOT U92 ( .A(n51), .Z(crcOut[18]) );
  GTECH_XOR3 U93 ( .A(crcIn[26]), .B(n52), .C(n53), .Z(n51) );
  GTECH_XOR3 U94 ( .A(crcIn[25]), .B(n43), .C(n53), .Z(crcOut[17]) );
  GTECH_XOR2 U95 ( .A(n40), .B(n33), .Z(n53) );
  GTECH_XOR2 U96 ( .A(n39), .B(n32), .Z(n33) );
  GTECH_XOR3 U97 ( .A(crcIn[24]), .B(n35), .C(n54), .Z(crcOut[16]) );
  GTECH_XOR3 U98 ( .A(crcIn[23]), .B(n28), .C(n35), .Z(crcOut[15]) );
  GTECH_XOR2 U99 ( .A(n37), .B(n43), .Z(n35) );
  GTECH_XOR2 U100 ( .A(crcIn[7]), .B(data[7]), .Z(n28) );
  GTECH_XOR3 U101 ( .A(crcIn[22]), .B(n30), .C(n52), .Z(crcOut[14]) );
  GTECH_XOR2 U102 ( .A(n37), .B(n49), .Z(n52) );
  GTECH_NOT U103 ( .A(n42), .Z(n49) );
  GTECH_XOR2 U104 ( .A(crcIn[6]), .B(data[6]), .Z(n42) );
  GTECH_NOT U105 ( .A(n44), .Z(n30) );
  GTECH_XOR3 U106 ( .A(crcIn[21]), .B(n32), .C(n40), .Z(crcOut[13]) );
  GTECH_XOR2 U107 ( .A(n41), .B(n44), .Z(n40) );
  GTECH_XOR2 U108 ( .A(crcIn[1]), .B(data[1]), .Z(n44) );
  GTECH_XOR2 U109 ( .A(crcIn[5]), .B(data[5]), .Z(n32) );
  GTECH_XOR2 U110 ( .A(crcIn[20]), .B(n54), .Z(crcOut[12]) );
  GTECH_XOR2 U111 ( .A(n39), .B(n41), .Z(n54) );
  GTECH_XOR2 U112 ( .A(crcIn[0]), .B(data[0]), .Z(n41) );
  GTECH_XOR2 U113 ( .A(crcIn[4]), .B(data[4]), .Z(n39) );
  GTECH_XOR2 U114 ( .A(crcIn[19]), .B(n43), .Z(crcOut[11]) );
  GTECH_XOR2 U115 ( .A(crcIn[3]), .B(data[3]), .Z(n43) );
  GTECH_XOR2 U116 ( .A(crcIn[18]), .B(n37), .Z(crcOut[10]) );
  GTECH_XOR2 U117 ( .A(crcIn[8]), .B(n37), .Z(crcOut[0]) );
  GTECH_XOR2 U118 ( .A(crcIn[2]), .B(data[2]), .Z(n37) );
endmodule

