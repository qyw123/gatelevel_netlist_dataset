
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_OAI21 U75 ( .A(n83), .B(n84), .C(n85), .Z(N155) );
  GTECH_OA22 U76 ( .A(n86), .B(n87), .C(n88), .D(n89), .Z(n85) );
  GTECH_NOT U77 ( .A(n90), .Z(n87) );
  GTECH_XOR2 U78 ( .A(n91), .B(n92), .Z(N154) );
  GTECH_NOT U79 ( .A(n83), .Z(n92) );
  GTECH_XOR2 U80 ( .A(n90), .B(n86), .Z(n83) );
  GTECH_AOI2N2 U81 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n86) );
  GTECH_NAND2 U82 ( .A(n95), .B(n96), .Z(n94) );
  GTECH_XOR2 U83 ( .A(n89), .B(n88), .Z(n90) );
  GTECH_AND2 U84 ( .A(n97), .B(n98), .Z(n88) );
  GTECH_OR_NOT U85 ( .A(n99), .B(n100), .Z(n98) );
  GTECH_OAI21 U86 ( .A(n101), .B(n100), .C(n102), .Z(n97) );
  GTECH_NAND2 U87 ( .A(I_b[7]), .B(I_a[7]), .Z(n89) );
  GTECH_NOT U88 ( .A(n84), .Z(n91) );
  GTECH_NAND2 U89 ( .A(n103), .B(n104), .Z(n84) );
  GTECH_XOR2 U90 ( .A(n104), .B(n103), .Z(N153) );
  GTECH_NOT U91 ( .A(n105), .Z(n103) );
  GTECH_XOR3 U92 ( .A(n106), .B(n95), .C(n93), .Z(n105) );
  GTECH_XOR3 U93 ( .A(n101), .B(n102), .C(n100), .Z(n93) );
  GTECH_OAI21 U94 ( .A(n107), .B(n108), .C(n109), .Z(n100) );
  GTECH_OAI21 U95 ( .A(n110), .B(n111), .C(n112), .Z(n109) );
  GTECH_NOT U96 ( .A(n111), .Z(n107) );
  GTECH_NOT U97 ( .A(n113), .Z(n102) );
  GTECH_NAND2 U98 ( .A(I_b[7]), .B(I_a[6]), .Z(n113) );
  GTECH_NOT U99 ( .A(n99), .Z(n101) );
  GTECH_NAND2 U100 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U101 ( .A(n114), .B(n115), .C(n116), .COUT(n95) );
  GTECH_NOT U102 ( .A(n117), .Z(n116) );
  GTECH_XOR2 U103 ( .A(n118), .B(n119), .Z(n115) );
  GTECH_AND2 U104 ( .A(I_a[7]), .B(I_b[5]), .Z(n119) );
  GTECH_NOT U105 ( .A(n96), .Z(n106) );
  GTECH_NAND2 U106 ( .A(I_a[7]), .B(n120), .Z(n96) );
  GTECH_NOT U107 ( .A(n121), .Z(n104) );
  GTECH_NAND2 U108 ( .A(n122), .B(n123), .Z(n121) );
  GTECH_NOT U109 ( .A(n124), .Z(n123) );
  GTECH_XOR2 U110 ( .A(n124), .B(n125), .Z(N152) );
  GTECH_NOT U111 ( .A(n122), .Z(n125) );
  GTECH_XOR4 U112 ( .A(n126), .B(n118), .C(n114), .D(n117), .Z(n122) );
  GTECH_XOR3 U113 ( .A(n110), .B(n112), .C(n111), .Z(n117) );
  GTECH_OAI21 U114 ( .A(n127), .B(n128), .C(n129), .Z(n111) );
  GTECH_OAI21 U115 ( .A(n130), .B(n131), .C(n132), .Z(n129) );
  GTECH_NOT U116 ( .A(n131), .Z(n127) );
  GTECH_NOT U117 ( .A(n133), .Z(n112) );
  GTECH_NAND2 U118 ( .A(I_b[7]), .B(I_a[5]), .Z(n133) );
  GTECH_NOT U119 ( .A(n108), .Z(n110) );
  GTECH_NAND2 U120 ( .A(I_b[6]), .B(I_a[6]), .Z(n108) );
  GTECH_ADD_ABC U121 ( .A(n134), .B(n135), .C(n136), .COUT(n114) );
  GTECH_NOT U122 ( .A(n137), .Z(n136) );
  GTECH_XOR3 U123 ( .A(n138), .B(n139), .C(n140), .Z(n135) );
  GTECH_NOT U124 ( .A(n120), .Z(n118) );
  GTECH_OAI21 U125 ( .A(n140), .B(n141), .C(n142), .Z(n120) );
  GTECH_OAI21 U126 ( .A(n138), .B(n143), .C(n139), .Z(n142) );
  GTECH_NOT U127 ( .A(n141), .Z(n138) );
  GTECH_NOT U128 ( .A(n143), .Z(n140) );
  GTECH_AND2 U129 ( .A(I_a[7]), .B(I_b[5]), .Z(n126) );
  GTECH_ADD_ABC U130 ( .A(n144), .B(n145), .C(n146), .COUT(n124) );
  GTECH_NOT U131 ( .A(n147), .Z(n146) );
  GTECH_OA22 U132 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n145) );
  GTECH_OA21 U133 ( .A(n152), .B(n153), .C(n154), .Z(n144) );
  GTECH_XOR3 U134 ( .A(n155), .B(n147), .C(n156), .Z(N151) );
  GTECH_OA21 U135 ( .A(n152), .B(n153), .C(n154), .Z(n156) );
  GTECH_OAI21 U136 ( .A(n157), .B(n158), .C(n159), .Z(n154) );
  GTECH_XOR2 U137 ( .A(n160), .B(n134), .Z(n147) );
  GTECH_ADD_ABC U138 ( .A(n161), .B(n162), .C(n163), .COUT(n134) );
  GTECH_NOT U139 ( .A(n164), .Z(n163) );
  GTECH_XOR3 U140 ( .A(n165), .B(n166), .C(n167), .Z(n162) );
  GTECH_XOR4 U141 ( .A(n139), .B(n143), .C(n141), .D(n137), .Z(n160) );
  GTECH_XOR3 U142 ( .A(n130), .B(n132), .C(n131), .Z(n137) );
  GTECH_OAI21 U143 ( .A(n168), .B(n169), .C(n170), .Z(n131) );
  GTECH_OAI21 U144 ( .A(n171), .B(n172), .C(n173), .Z(n170) );
  GTECH_NOT U145 ( .A(n172), .Z(n168) );
  GTECH_NOT U146 ( .A(n174), .Z(n132) );
  GTECH_NAND2 U147 ( .A(I_b[7]), .B(I_a[4]), .Z(n174) );
  GTECH_NOT U148 ( .A(n128), .Z(n130) );
  GTECH_NAND2 U149 ( .A(I_b[6]), .B(I_a[5]), .Z(n128) );
  GTECH_NAND2 U150 ( .A(I_a[7]), .B(I_b[4]), .Z(n141) );
  GTECH_OAI21 U151 ( .A(n167), .B(n175), .C(n176), .Z(n143) );
  GTECH_OAI21 U152 ( .A(n165), .B(n177), .C(n166), .Z(n176) );
  GTECH_NOT U153 ( .A(n175), .Z(n165) );
  GTECH_NOT U154 ( .A(n177), .Z(n167) );
  GTECH_NOT U155 ( .A(n178), .Z(n139) );
  GTECH_NAND2 U156 ( .A(I_a[6]), .B(I_b[5]), .Z(n178) );
  GTECH_OA22 U157 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n155) );
  GTECH_NOT U158 ( .A(n179), .Z(n151) );
  GTECH_NOT U159 ( .A(I_a[7]), .Z(n149) );
  GTECH_XOR3 U160 ( .A(n152), .B(n157), .C(n180), .Z(N150) );
  GTECH_NOT U161 ( .A(n159), .Z(n180) );
  GTECH_XOR2 U162 ( .A(n181), .B(n161), .Z(n159) );
  GTECH_ADD_ABC U163 ( .A(n182), .B(n183), .C(n184), .COUT(n161) );
  GTECH_NOT U164 ( .A(n185), .Z(n184) );
  GTECH_XOR3 U165 ( .A(n186), .B(n187), .C(n188), .Z(n183) );
  GTECH_XOR4 U166 ( .A(n166), .B(n177), .C(n175), .D(n164), .Z(n181) );
  GTECH_XOR3 U167 ( .A(n171), .B(n173), .C(n172), .Z(n164) );
  GTECH_OAI21 U168 ( .A(n189), .B(n190), .C(n191), .Z(n172) );
  GTECH_OAI21 U169 ( .A(n192), .B(n193), .C(n194), .Z(n191) );
  GTECH_NOT U170 ( .A(n193), .Z(n189) );
  GTECH_NOT U171 ( .A(n195), .Z(n173) );
  GTECH_NAND2 U172 ( .A(I_b[7]), .B(I_a[3]), .Z(n195) );
  GTECH_NOT U173 ( .A(n169), .Z(n171) );
  GTECH_NAND2 U174 ( .A(I_b[6]), .B(I_a[4]), .Z(n169) );
  GTECH_NAND2 U175 ( .A(I_a[6]), .B(I_b[4]), .Z(n175) );
  GTECH_OAI21 U176 ( .A(n188), .B(n196), .C(n197), .Z(n177) );
  GTECH_OAI21 U177 ( .A(n186), .B(n198), .C(n187), .Z(n197) );
  GTECH_NOT U178 ( .A(n196), .Z(n186) );
  GTECH_NOT U179 ( .A(n198), .Z(n188) );
  GTECH_NOT U180 ( .A(n199), .Z(n166) );
  GTECH_NAND2 U181 ( .A(I_a[5]), .B(I_b[5]), .Z(n199) );
  GTECH_NOT U182 ( .A(n153), .Z(n157) );
  GTECH_XOR2 U183 ( .A(n179), .B(n150), .Z(n153) );
  GTECH_AOI2N2 U184 ( .A(n200), .B(n201), .C(n202), .D(n203), .Z(n150) );
  GTECH_NAND2 U185 ( .A(n202), .B(n203), .Z(n201) );
  GTECH_XOR2 U186 ( .A(n204), .B(n148), .Z(n179) );
  GTECH_AND2 U187 ( .A(n205), .B(n206), .Z(n148) );
  GTECH_OR_NOT U188 ( .A(n207), .B(n208), .Z(n206) );
  GTECH_OAI21 U189 ( .A(n209), .B(n208), .C(n210), .Z(n205) );
  GTECH_NAND2 U190 ( .A(I_a[7]), .B(I_b[3]), .Z(n204) );
  GTECH_NOT U191 ( .A(n158), .Z(n152) );
  GTECH_OAI2N2 U192 ( .A(n211), .B(n212), .C(n213), .D(n214), .Z(n158) );
  GTECH_NAND2 U193 ( .A(n211), .B(n212), .Z(n214) );
  GTECH_XOR3 U194 ( .A(n211), .B(n215), .C(n216), .Z(N149) );
  GTECH_NOT U195 ( .A(n213), .Z(n216) );
  GTECH_XOR2 U196 ( .A(n217), .B(n182), .Z(n213) );
  GTECH_ADD_ABC U197 ( .A(n218), .B(n219), .C(n220), .COUT(n182) );
  GTECH_XOR3 U198 ( .A(n221), .B(n222), .C(n223), .Z(n219) );
  GTECH_OA21 U199 ( .A(n224), .B(n225), .C(n226), .Z(n218) );
  GTECH_XOR4 U200 ( .A(n187), .B(n198), .C(n196), .D(n185), .Z(n217) );
  GTECH_XOR3 U201 ( .A(n192), .B(n194), .C(n193), .Z(n185) );
  GTECH_OAI21 U202 ( .A(n227), .B(n228), .C(n229), .Z(n193) );
  GTECH_NOT U203 ( .A(n230), .Z(n194) );
  GTECH_NAND2 U204 ( .A(I_b[7]), .B(I_a[2]), .Z(n230) );
  GTECH_NOT U205 ( .A(n190), .Z(n192) );
  GTECH_NAND2 U206 ( .A(I_b[6]), .B(I_a[3]), .Z(n190) );
  GTECH_NAND2 U207 ( .A(I_a[5]), .B(I_b[4]), .Z(n196) );
  GTECH_OAI21 U208 ( .A(n223), .B(n231), .C(n232), .Z(n198) );
  GTECH_OAI21 U209 ( .A(n221), .B(n233), .C(n222), .Z(n232) );
  GTECH_NOT U210 ( .A(n231), .Z(n221) );
  GTECH_NOT U211 ( .A(n233), .Z(n223) );
  GTECH_NOT U212 ( .A(n234), .Z(n187) );
  GTECH_NAND2 U213 ( .A(I_b[5]), .B(I_a[4]), .Z(n234) );
  GTECH_NOT U214 ( .A(n212), .Z(n215) );
  GTECH_XOR3 U215 ( .A(n235), .B(n202), .C(n200), .Z(n212) );
  GTECH_XOR3 U216 ( .A(n209), .B(n210), .C(n208), .Z(n200) );
  GTECH_OAI21 U217 ( .A(n236), .B(n237), .C(n238), .Z(n208) );
  GTECH_OAI21 U218 ( .A(n239), .B(n240), .C(n241), .Z(n238) );
  GTECH_NOT U219 ( .A(n240), .Z(n236) );
  GTECH_NOT U220 ( .A(n242), .Z(n210) );
  GTECH_NAND2 U221 ( .A(I_a[6]), .B(I_b[3]), .Z(n242) );
  GTECH_NOT U222 ( .A(n207), .Z(n209) );
  GTECH_NAND2 U223 ( .A(I_a[7]), .B(I_b[2]), .Z(n207) );
  GTECH_ADD_ABC U224 ( .A(n243), .B(n244), .C(n245), .COUT(n202) );
  GTECH_XOR2 U225 ( .A(n246), .B(n247), .Z(n244) );
  GTECH_AND2 U226 ( .A(I_a[7]), .B(I_b[1]), .Z(n247) );
  GTECH_NOT U227 ( .A(n203), .Z(n235) );
  GTECH_NAND2 U228 ( .A(I_a[7]), .B(n248), .Z(n203) );
  GTECH_ADD_ABC U229 ( .A(n249), .B(n250), .C(n251), .COUT(n211) );
  GTECH_XOR3 U230 ( .A(n243), .B(n252), .C(n245), .Z(n250) );
  GTECH_NOT U231 ( .A(n253), .Z(n245) );
  GTECH_XOR2 U232 ( .A(n249), .B(n254), .Z(N148) );
  GTECH_XOR4 U233 ( .A(n252), .B(n253), .C(n251), .D(n243), .Z(n254) );
  GTECH_ADD_ABC U234 ( .A(n255), .B(n256), .C(n257), .COUT(n243) );
  GTECH_XOR3 U235 ( .A(n258), .B(n259), .C(n260), .Z(n256) );
  GTECH_XOR2 U236 ( .A(n261), .B(n262), .Z(n251) );
  GTECH_OA21 U237 ( .A(n224), .B(n225), .C(n226), .Z(n262) );
  GTECH_OAI21 U238 ( .A(n263), .B(n264), .C(n265), .Z(n226) );
  GTECH_NOT U239 ( .A(n224), .Z(n264) );
  GTECH_XOR4 U240 ( .A(n222), .B(n233), .C(n231), .D(n220), .Z(n261) );
  GTECH_XOR3 U241 ( .A(n266), .B(n267), .C(n229), .Z(n220) );
  GTECH_NAND3 U242 ( .A(I_b[6]), .B(I_a[1]), .C(n268), .Z(n229) );
  GTECH_NOT U243 ( .A(n228), .Z(n267) );
  GTECH_NAND2 U244 ( .A(I_b[7]), .B(I_a[1]), .Z(n228) );
  GTECH_NOT U245 ( .A(n227), .Z(n266) );
  GTECH_NAND2 U246 ( .A(I_b[6]), .B(I_a[2]), .Z(n227) );
  GTECH_NAND2 U247 ( .A(I_b[4]), .B(I_a[4]), .Z(n231) );
  GTECH_OAI21 U248 ( .A(n269), .B(n270), .C(n271), .Z(n233) );
  GTECH_OAI21 U249 ( .A(n272), .B(n273), .C(n274), .Z(n271) );
  GTECH_NOT U250 ( .A(n273), .Z(n269) );
  GTECH_NOT U251 ( .A(n275), .Z(n222) );
  GTECH_NAND2 U252 ( .A(I_b[5]), .B(I_a[3]), .Z(n275) );
  GTECH_XOR3 U253 ( .A(n239), .B(n241), .C(n240), .Z(n253) );
  GTECH_OAI21 U254 ( .A(n276), .B(n277), .C(n278), .Z(n240) );
  GTECH_OAI21 U255 ( .A(n279), .B(n280), .C(n281), .Z(n278) );
  GTECH_NOT U256 ( .A(n280), .Z(n276) );
  GTECH_NOT U257 ( .A(n282), .Z(n241) );
  GTECH_NAND2 U258 ( .A(I_a[5]), .B(I_b[3]), .Z(n282) );
  GTECH_NOT U259 ( .A(n237), .Z(n239) );
  GTECH_NAND2 U260 ( .A(I_a[6]), .B(I_b[2]), .Z(n237) );
  GTECH_XOR2 U261 ( .A(n283), .B(n246), .Z(n252) );
  GTECH_NOT U262 ( .A(n248), .Z(n246) );
  GTECH_OAI21 U263 ( .A(n260), .B(n284), .C(n285), .Z(n248) );
  GTECH_OAI21 U264 ( .A(n258), .B(n286), .C(n259), .Z(n285) );
  GTECH_NOT U265 ( .A(n286), .Z(n260) );
  GTECH_AND2 U266 ( .A(I_a[7]), .B(I_b[1]), .Z(n283) );
  GTECH_ADD_ABC U267 ( .A(n287), .B(n288), .C(n289), .COUT(n249) );
  GTECH_NOT U268 ( .A(n290), .Z(n289) );
  GTECH_XOR3 U269 ( .A(n255), .B(n291), .C(n257), .Z(n288) );
  GTECH_NOT U270 ( .A(n292), .Z(n257) );
  GTECH_NOT U271 ( .A(n293), .Z(n291) );
  GTECH_XOR2 U272 ( .A(n294), .B(n287), .Z(N147) );
  GTECH_ADD_ABC U273 ( .A(n295), .B(n296), .C(n297), .COUT(n287) );
  GTECH_XOR3 U274 ( .A(n298), .B(n299), .C(n300), .Z(n296) );
  GTECH_OA21 U275 ( .A(n301), .B(n302), .C(n303), .Z(n295) );
  GTECH_XOR4 U276 ( .A(n292), .B(n255), .C(n293), .D(n290), .Z(n294) );
  GTECH_XOR3 U277 ( .A(n265), .B(n225), .C(n224), .Z(n290) );
  GTECH_XOR2 U278 ( .A(n304), .B(n268), .Z(n224) );
  GTECH_NOT U279 ( .A(n305), .Z(n268) );
  GTECH_NAND2 U280 ( .A(I_b[7]), .B(I_a[0]), .Z(n305) );
  GTECH_NAND2 U281 ( .A(I_b[6]), .B(I_a[1]), .Z(n304) );
  GTECH_NOT U282 ( .A(n263), .Z(n225) );
  GTECH_XOR3 U283 ( .A(n272), .B(n274), .C(n273), .Z(n263) );
  GTECH_OAI21 U284 ( .A(n306), .B(n307), .C(n308), .Z(n273) );
  GTECH_NOT U285 ( .A(n309), .Z(n274) );
  GTECH_NAND2 U286 ( .A(I_b[5]), .B(I_a[2]), .Z(n309) );
  GTECH_NOT U287 ( .A(n270), .Z(n272) );
  GTECH_NAND2 U288 ( .A(I_b[4]), .B(I_a[3]), .Z(n270) );
  GTECH_NOT U289 ( .A(n310), .Z(n265) );
  GTECH_NAND3 U290 ( .A(I_a[0]), .B(n311), .C(I_b[6]), .Z(n310) );
  GTECH_NOT U291 ( .A(n312), .Z(n311) );
  GTECH_XOR3 U292 ( .A(n258), .B(n259), .C(n286), .Z(n293) );
  GTECH_OAI21 U293 ( .A(n313), .B(n314), .C(n315), .Z(n286) );
  GTECH_OAI21 U294 ( .A(n316), .B(n317), .C(n318), .Z(n315) );
  GTECH_NOT U295 ( .A(n319), .Z(n259) );
  GTECH_NAND2 U296 ( .A(I_a[6]), .B(I_b[1]), .Z(n319) );
  GTECH_NOT U297 ( .A(n284), .Z(n258) );
  GTECH_NAND2 U298 ( .A(I_a[7]), .B(I_b[0]), .Z(n284) );
  GTECH_ADD_ABC U299 ( .A(n298), .B(n320), .C(n300), .COUT(n255) );
  GTECH_NOT U300 ( .A(n321), .Z(n300) );
  GTECH_XOR3 U301 ( .A(n316), .B(n318), .C(n313), .Z(n320) );
  GTECH_NOT U302 ( .A(n317), .Z(n313) );
  GTECH_XOR3 U303 ( .A(n279), .B(n281), .C(n280), .Z(n292) );
  GTECH_OAI21 U304 ( .A(n322), .B(n323), .C(n324), .Z(n280) );
  GTECH_OAI21 U305 ( .A(n325), .B(n326), .C(n327), .Z(n324) );
  GTECH_NOT U306 ( .A(n326), .Z(n322) );
  GTECH_NOT U307 ( .A(n328), .Z(n281) );
  GTECH_NAND2 U308 ( .A(I_b[3]), .B(I_a[4]), .Z(n328) );
  GTECH_NOT U309 ( .A(n277), .Z(n279) );
  GTECH_NAND2 U310 ( .A(I_a[5]), .B(I_b[2]), .Z(n277) );
  GTECH_XOR2 U311 ( .A(n329), .B(n330), .Z(N146) );
  GTECH_XOR4 U312 ( .A(n299), .B(n321), .C(n297), .D(n298), .Z(n330) );
  GTECH_ADD_ABC U313 ( .A(n331), .B(n332), .C(n333), .COUT(n298) );
  GTECH_NOT U314 ( .A(n334), .Z(n333) );
  GTECH_XOR3 U315 ( .A(n335), .B(n336), .C(n337), .Z(n332) );
  GTECH_XOR2 U316 ( .A(n312), .B(n338), .Z(n297) );
  GTECH_AND2 U317 ( .A(I_b[6]), .B(I_a[0]), .Z(n338) );
  GTECH_XOR3 U318 ( .A(n339), .B(n340), .C(n308), .Z(n312) );
  GTECH_NAND3 U319 ( .A(I_b[4]), .B(I_a[1]), .C(n341), .Z(n308) );
  GTECH_NOT U320 ( .A(n307), .Z(n340) );
  GTECH_NAND2 U321 ( .A(I_b[5]), .B(I_a[1]), .Z(n307) );
  GTECH_NOT U322 ( .A(n306), .Z(n339) );
  GTECH_NAND2 U323 ( .A(I_b[4]), .B(I_a[2]), .Z(n306) );
  GTECH_XOR3 U324 ( .A(n325), .B(n327), .C(n326), .Z(n321) );
  GTECH_OAI21 U325 ( .A(n342), .B(n343), .C(n344), .Z(n326) );
  GTECH_OAI21 U326 ( .A(n345), .B(n346), .C(n347), .Z(n344) );
  GTECH_NOT U327 ( .A(n346), .Z(n342) );
  GTECH_NOT U328 ( .A(n348), .Z(n327) );
  GTECH_NAND2 U329 ( .A(I_b[3]), .B(I_a[3]), .Z(n348) );
  GTECH_NOT U330 ( .A(n323), .Z(n325) );
  GTECH_NAND2 U331 ( .A(I_b[2]), .B(I_a[4]), .Z(n323) );
  GTECH_NOT U332 ( .A(n349), .Z(n299) );
  GTECH_XOR3 U333 ( .A(n316), .B(n318), .C(n317), .Z(n349) );
  GTECH_OAI21 U334 ( .A(n337), .B(n350), .C(n351), .Z(n317) );
  GTECH_OAI21 U335 ( .A(n335), .B(n352), .C(n336), .Z(n351) );
  GTECH_NOT U336 ( .A(n350), .Z(n335) );
  GTECH_NOT U337 ( .A(n352), .Z(n337) );
  GTECH_NOT U338 ( .A(n353), .Z(n318) );
  GTECH_NAND2 U339 ( .A(I_a[5]), .B(I_b[1]), .Z(n353) );
  GTECH_NOT U340 ( .A(n314), .Z(n316) );
  GTECH_NAND2 U341 ( .A(I_a[6]), .B(I_b[0]), .Z(n314) );
  GTECH_OA21 U342 ( .A(n301), .B(n302), .C(n303), .Z(n329) );
  GTECH_OAI21 U343 ( .A(n354), .B(n355), .C(n356), .Z(n303) );
  GTECH_NOT U344 ( .A(n301), .Z(n355) );
  GTECH_XOR3 U345 ( .A(n356), .B(n302), .C(n301), .Z(N145) );
  GTECH_XOR2 U346 ( .A(n357), .B(n341), .Z(n301) );
  GTECH_NOT U347 ( .A(n358), .Z(n341) );
  GTECH_NAND2 U348 ( .A(I_b[5]), .B(I_a[0]), .Z(n358) );
  GTECH_NAND2 U349 ( .A(I_b[4]), .B(I_a[1]), .Z(n357) );
  GTECH_NOT U350 ( .A(n354), .Z(n302) );
  GTECH_XOR2 U351 ( .A(n359), .B(n331), .Z(n354) );
  GTECH_ADD_ABC U352 ( .A(n360), .B(n361), .C(n362), .COUT(n331) );
  GTECH_XOR3 U353 ( .A(n363), .B(n364), .C(n365), .Z(n361) );
  GTECH_OA21 U354 ( .A(n366), .B(n367), .C(n368), .Z(n360) );
  GTECH_XOR4 U355 ( .A(n336), .B(n352), .C(n350), .D(n334), .Z(n359) );
  GTECH_XOR3 U356 ( .A(n345), .B(n347), .C(n346), .Z(n334) );
  GTECH_OAI21 U357 ( .A(n369), .B(n370), .C(n371), .Z(n346) );
  GTECH_NOT U358 ( .A(n372), .Z(n347) );
  GTECH_NAND2 U359 ( .A(I_b[3]), .B(I_a[2]), .Z(n372) );
  GTECH_NOT U360 ( .A(n343), .Z(n345) );
  GTECH_NAND2 U361 ( .A(I_b[2]), .B(I_a[3]), .Z(n343) );
  GTECH_NAND2 U362 ( .A(I_a[5]), .B(I_b[0]), .Z(n350) );
  GTECH_OAI21 U363 ( .A(n365), .B(n373), .C(n374), .Z(n352) );
  GTECH_OAI21 U364 ( .A(n363), .B(n375), .C(n364), .Z(n374) );
  GTECH_NOT U365 ( .A(n375), .Z(n365) );
  GTECH_NOT U366 ( .A(n376), .Z(n336) );
  GTECH_NAND2 U367 ( .A(I_a[4]), .B(I_b[1]), .Z(n376) );
  GTECH_NOT U368 ( .A(n377), .Z(n356) );
  GTECH_NAND3 U369 ( .A(I_a[0]), .B(n378), .C(I_b[4]), .Z(n377) );
  GTECH_XOR2 U370 ( .A(n379), .B(n378), .Z(N144) );
  GTECH_XOR2 U371 ( .A(n380), .B(n381), .Z(n378) );
  GTECH_XOR4 U372 ( .A(n364), .B(n375), .C(n362), .D(n363), .Z(n381) );
  GTECH_NOT U373 ( .A(n373), .Z(n363) );
  GTECH_NAND2 U374 ( .A(I_a[4]), .B(I_b[0]), .Z(n373) );
  GTECH_XOR3 U375 ( .A(n382), .B(n383), .C(n371), .Z(n362) );
  GTECH_NAND3 U376 ( .A(I_b[2]), .B(I_a[1]), .C(n384), .Z(n371) );
  GTECH_NOT U377 ( .A(n370), .Z(n383) );
  GTECH_NAND2 U378 ( .A(I_b[3]), .B(I_a[1]), .Z(n370) );
  GTECH_NOT U379 ( .A(n369), .Z(n382) );
  GTECH_NAND2 U380 ( .A(I_b[2]), .B(I_a[2]), .Z(n369) );
  GTECH_OAI21 U381 ( .A(n385), .B(n386), .C(n387), .Z(n375) );
  GTECH_OAI21 U382 ( .A(n388), .B(n389), .C(n390), .Z(n387) );
  GTECH_NOT U383 ( .A(n389), .Z(n385) );
  GTECH_NOT U384 ( .A(n391), .Z(n364) );
  GTECH_NAND2 U385 ( .A(I_a[3]), .B(I_b[1]), .Z(n391) );
  GTECH_OA21 U386 ( .A(n366), .B(n367), .C(n368), .Z(n380) );
  GTECH_OAI21 U387 ( .A(n392), .B(n393), .C(n394), .Z(n368) );
  GTECH_NOT U388 ( .A(n366), .Z(n393) );
  GTECH_AND2 U389 ( .A(I_b[4]), .B(I_a[0]), .Z(n379) );
  GTECH_XOR3 U390 ( .A(n394), .B(n367), .C(n366), .Z(N143) );
  GTECH_XOR2 U391 ( .A(n395), .B(n384), .Z(n366) );
  GTECH_NOT U392 ( .A(n396), .Z(n384) );
  GTECH_NAND2 U393 ( .A(I_b[3]), .B(I_a[0]), .Z(n396) );
  GTECH_NAND2 U394 ( .A(I_b[2]), .B(I_a[1]), .Z(n395) );
  GTECH_NOT U395 ( .A(n392), .Z(n367) );
  GTECH_XOR3 U396 ( .A(n388), .B(n390), .C(n389), .Z(n392) );
  GTECH_OAI21 U397 ( .A(n397), .B(n398), .C(n399), .Z(n389) );
  GTECH_NOT U398 ( .A(n400), .Z(n390) );
  GTECH_NAND2 U399 ( .A(I_b[1]), .B(I_a[2]), .Z(n400) );
  GTECH_NOT U400 ( .A(n386), .Z(n388) );
  GTECH_NAND2 U401 ( .A(I_b[0]), .B(I_a[3]), .Z(n386) );
  GTECH_NOT U402 ( .A(n401), .Z(n394) );
  GTECH_NAND3 U403 ( .A(I_a[0]), .B(n402), .C(I_b[2]), .Z(n401) );
  GTECH_XOR2 U404 ( .A(n403), .B(n402), .Z(N142) );
  GTECH_NOT U405 ( .A(n404), .Z(n402) );
  GTECH_XOR3 U406 ( .A(n405), .B(n406), .C(n399), .Z(n404) );
  GTECH_NAND3 U407 ( .A(n407), .B(I_b[0]), .C(I_a[1]), .Z(n399) );
  GTECH_NOT U408 ( .A(n397), .Z(n406) );
  GTECH_NAND2 U409 ( .A(I_a[1]), .B(I_b[1]), .Z(n397) );
  GTECH_NOT U410 ( .A(n398), .Z(n405) );
  GTECH_NAND2 U411 ( .A(I_b[0]), .B(I_a[2]), .Z(n398) );
  GTECH_AND2 U412 ( .A(I_b[2]), .B(I_a[0]), .Z(n403) );
  GTECH_XOR2 U413 ( .A(n407), .B(n408), .Z(N141) );
  GTECH_AND2 U414 ( .A(I_a[1]), .B(I_b[0]), .Z(n408) );
  GTECH_NOT U415 ( .A(n409), .Z(n407) );
  GTECH_NAND2 U416 ( .A(I_a[0]), .B(I_b[1]), .Z(n409) );
  GTECH_AND2 U417 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

