
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378;

  GTECH_MUX2 U133 ( .A(n272), .B(n273), .S(n274), .Z(sum[9]) );
  GTECH_XNOR2 U134 ( .A(n275), .B(n276), .Z(n273) );
  GTECH_XOR2 U135 ( .A(n275), .B(n277), .Z(n272) );
  GTECH_NOR2 U136 ( .A(n278), .B(n279), .Z(n275) );
  GTECH_NAND2 U137 ( .A(n280), .B(n281), .Z(sum[8]) );
  GTECH_AO21 U138 ( .A(n276), .B(n277), .C(n274), .Z(n280) );
  GTECH_MUX2 U139 ( .A(n282), .B(n283), .S(n284), .Z(sum[7]) );
  GTECH_XOR2 U140 ( .A(n285), .B(n286), .Z(n283) );
  GTECH_XOR2 U141 ( .A(n287), .B(n285), .Z(n282) );
  GTECH_XOR2 U142 ( .A(a[7]), .B(b[7]), .Z(n285) );
  GTECH_OA21 U143 ( .A(a[6]), .B(n288), .C(n289), .Z(n287) );
  GTECH_AO21 U144 ( .A(n288), .B(a[6]), .C(b[6]), .Z(n289) );
  GTECH_MUX2 U145 ( .A(n290), .B(n291), .S(n284), .Z(sum[6]) );
  GTECH_XOR2 U146 ( .A(n292), .B(n293), .Z(n291) );
  GTECH_XNOR2 U147 ( .A(n292), .B(n288), .Z(n290) );
  GTECH_OAI21 U148 ( .A(n294), .B(n295), .C(n296), .Z(n288) );
  GTECH_XOR2 U149 ( .A(a[6]), .B(n297), .Z(n292) );
  GTECH_MUX2 U150 ( .A(n298), .B(n299), .S(n300), .Z(sum[5]) );
  GTECH_AND_NOT U151 ( .A(n296), .B(n294), .Z(n300) );
  GTECH_OAI21 U152 ( .A(n301), .B(n284), .C(n302), .Z(n299) );
  GTECH_OAI21 U153 ( .A(n303), .B(n304), .C(n295), .Z(n298) );
  GTECH_XNOR2 U154 ( .A(n305), .B(n284), .Z(sum[4]) );
  GTECH_MUX2 U155 ( .A(n306), .B(n307), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U156 ( .A(n308), .B(n309), .Z(n307) );
  GTECH_XOR2 U157 ( .A(n308), .B(n310), .Z(n306) );
  GTECH_OA21 U158 ( .A(n311), .B(n312), .C(n313), .Z(n310) );
  GTECH_XNOR2 U159 ( .A(a[3]), .B(b[3]), .Z(n308) );
  GTECH_MUX2 U160 ( .A(n314), .B(n315), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U161 ( .A(n316), .B(n317), .Z(n315) );
  GTECH_XNOR2 U162 ( .A(n312), .B(n317), .Z(n314) );
  GTECH_AND_NOT U163 ( .A(n313), .B(n311), .Z(n317) );
  GTECH_OA21 U164 ( .A(n318), .B(n319), .C(n320), .Z(n312) );
  GTECH_MUX2 U165 ( .A(n321), .B(n322), .S(n323), .Z(sum[1]) );
  GTECH_AND_NOT U166 ( .A(n320), .B(n318), .Z(n323) );
  GTECH_AO21 U167 ( .A(n324), .B(n319), .C(n325), .Z(n322) );
  GTECH_OAI21 U168 ( .A(n325), .B(n324), .C(n319), .Z(n321) );
  GTECH_NAND2 U169 ( .A(a[0]), .B(b[0]), .Z(n319) );
  GTECH_NOT U170 ( .A(cin), .Z(n324) );
  GTECH_MUX2 U171 ( .A(n326), .B(n327), .S(n328), .Z(sum[15]) );
  GTECH_XOR2 U172 ( .A(n329), .B(n330), .Z(n327) );
  GTECH_AOI21 U173 ( .A(n331), .B(n332), .C(n333), .Z(n330) );
  GTECH_XNOR2 U174 ( .A(n329), .B(n334), .Z(n326) );
  GTECH_XNOR2 U175 ( .A(a[15]), .B(b[15]), .Z(n329) );
  GTECH_MUX2 U176 ( .A(n335), .B(n336), .S(n328), .Z(sum[14]) );
  GTECH_XOR2 U177 ( .A(n337), .B(n332), .Z(n336) );
  GTECH_AOI21 U178 ( .A(n338), .B(n339), .C(n340), .Z(n332) );
  GTECH_XOR2 U179 ( .A(n337), .B(n341), .Z(n335) );
  GTECH_NOR2 U180 ( .A(n342), .B(n333), .Z(n337) );
  GTECH_MUX2 U181 ( .A(n343), .B(n344), .S(n328), .Z(sum[13]) );
  GTECH_XOR2 U182 ( .A(n345), .B(n339), .Z(n344) );
  GTECH_XNOR2 U183 ( .A(n345), .B(n346), .Z(n343) );
  GTECH_OAI21 U184 ( .A(a[13]), .B(b[13]), .C(n338), .Z(n345) );
  GTECH_NAND2 U185 ( .A(n347), .B(n348), .Z(sum[12]) );
  GTECH_AO21 U186 ( .A(n339), .B(n346), .C(n328), .Z(n347) );
  GTECH_MUX2 U187 ( .A(n349), .B(n350), .S(n274), .Z(sum[11]) );
  GTECH_XOR2 U188 ( .A(n351), .B(n352), .Z(n350) );
  GTECH_AOI21 U189 ( .A(n353), .B(n354), .C(n355), .Z(n352) );
  GTECH_XNOR2 U190 ( .A(n351), .B(n356), .Z(n349) );
  GTECH_XNOR2 U191 ( .A(a[11]), .B(b[11]), .Z(n351) );
  GTECH_MUX2 U192 ( .A(n357), .B(n358), .S(n274), .Z(sum[10]) );
  GTECH_XOR2 U193 ( .A(n354), .B(n359), .Z(n358) );
  GTECH_AO21 U194 ( .A(n360), .B(n361), .C(n279), .Z(n354) );
  GTECH_XOR2 U195 ( .A(n362), .B(n359), .Z(n357) );
  GTECH_NOR2 U196 ( .A(n363), .B(n355), .Z(n359) );
  GTECH_XNOR2 U197 ( .A(cin), .B(n364), .Z(sum[0]) );
  GTECH_OAI21 U198 ( .A(n328), .B(n365), .C(n348), .Z(cout) );
  GTECH_NAND3 U199 ( .A(n339), .B(n346), .C(n328), .Z(n348) );
  GTECH_NOT U200 ( .A(n366), .Z(n346) );
  GTECH_NAND2 U201 ( .A(a[12]), .B(b[12]), .Z(n339) );
  GTECH_AOI21 U202 ( .A(n334), .B(a[15]), .C(n367), .Z(n365) );
  GTECH_OA21 U203 ( .A(a[15]), .B(n334), .C(b[15]), .Z(n367) );
  GTECH_AO21 U204 ( .A(n331), .B(n341), .C(n333), .Z(n334) );
  GTECH_AND2 U205 ( .A(a[14]), .B(b[14]), .Z(n333) );
  GTECH_AOI21 U206 ( .A(n338), .B(n366), .C(n340), .Z(n341) );
  GTECH_NOR2 U207 ( .A(b[13]), .B(a[13]), .Z(n340) );
  GTECH_NOR2 U208 ( .A(b[12]), .B(a[12]), .Z(n366) );
  GTECH_NAND2 U209 ( .A(a[13]), .B(b[13]), .Z(n338) );
  GTECH_NOT U210 ( .A(n342), .Z(n331) );
  GTECH_NOR2 U211 ( .A(a[14]), .B(b[14]), .Z(n342) );
  GTECH_OA21 U212 ( .A(n368), .B(n274), .C(n281), .Z(n328) );
  GTECH_NAND3 U213 ( .A(n276), .B(n277), .C(n274), .Z(n281) );
  GTECH_NOT U214 ( .A(n361), .Z(n276) );
  GTECH_AND2 U215 ( .A(b[8]), .B(a[8]), .Z(n361) );
  GTECH_MUX2 U216 ( .A(n305), .B(n369), .S(n284), .Z(n274) );
  GTECH_NOT U217 ( .A(n304), .Z(n284) );
  GTECH_MUX2 U218 ( .A(n364), .B(n370), .S(cin), .Z(n304) );
  GTECH_AOI21 U219 ( .A(n309), .B(a[3]), .C(n371), .Z(n370) );
  GTECH_OA21 U220 ( .A(a[3]), .B(n309), .C(b[3]), .Z(n371) );
  GTECH_OAI21 U221 ( .A(n316), .B(n311), .C(n313), .Z(n309) );
  GTECH_NAND2 U222 ( .A(a[2]), .B(b[2]), .Z(n313) );
  GTECH_NOR2 U223 ( .A(a[2]), .B(b[2]), .Z(n311) );
  GTECH_OA21 U224 ( .A(n318), .B(n325), .C(n320), .Z(n316) );
  GTECH_NAND2 U225 ( .A(a[1]), .B(b[1]), .Z(n320) );
  GTECH_AND_NOT U226 ( .A(n372), .B(a[0]), .Z(n325) );
  GTECH_NOR2 U227 ( .A(a[1]), .B(b[1]), .Z(n318) );
  GTECH_XNOR2 U228 ( .A(n373), .B(n372), .Z(n364) );
  GTECH_NOT U229 ( .A(b[0]), .Z(n372) );
  GTECH_NOT U230 ( .A(a[0]), .Z(n373) );
  GTECH_AOI21 U231 ( .A(n286), .B(a[7]), .C(n374), .Z(n369) );
  GTECH_OA21 U232 ( .A(a[7]), .B(n286), .C(b[7]), .Z(n374) );
  GTECH_OAI21 U233 ( .A(n293), .B(n375), .C(n376), .Z(n286) );
  GTECH_AO21 U234 ( .A(n375), .B(n293), .C(n297), .Z(n376) );
  GTECH_NOT U235 ( .A(b[6]), .Z(n297) );
  GTECH_NOT U236 ( .A(a[6]), .Z(n375) );
  GTECH_OA21 U237 ( .A(n303), .B(n294), .C(n296), .Z(n293) );
  GTECH_NAND2 U238 ( .A(a[5]), .B(b[5]), .Z(n296) );
  GTECH_NOR2 U239 ( .A(a[5]), .B(b[5]), .Z(n294) );
  GTECH_NAND2 U240 ( .A(n295), .B(n302), .Z(n305) );
  GTECH_NOT U241 ( .A(n303), .Z(n302) );
  GTECH_NOR2 U242 ( .A(a[4]), .B(b[4]), .Z(n303) );
  GTECH_NOT U243 ( .A(n301), .Z(n295) );
  GTECH_AND2 U244 ( .A(a[4]), .B(b[4]), .Z(n301) );
  GTECH_AOI21 U245 ( .A(n356), .B(a[11]), .C(n377), .Z(n368) );
  GTECH_OA21 U246 ( .A(a[11]), .B(n356), .C(b[11]), .Z(n377) );
  GTECH_AO21 U247 ( .A(n362), .B(n353), .C(n355), .Z(n356) );
  GTECH_AND2 U248 ( .A(a[10]), .B(b[10]), .Z(n355) );
  GTECH_NOT U249 ( .A(n363), .Z(n353) );
  GTECH_NOR2 U250 ( .A(a[10]), .B(b[10]), .Z(n363) );
  GTECH_AO21 U251 ( .A(n277), .B(n360), .C(n279), .Z(n362) );
  GTECH_AND2 U252 ( .A(a[9]), .B(b[9]), .Z(n279) );
  GTECH_NOT U253 ( .A(n278), .Z(n360) );
  GTECH_NOR2 U254 ( .A(a[9]), .B(b[9]), .Z(n278) );
  GTECH_OR_NOT U255 ( .A(b[8]), .B(n378), .Z(n277) );
  GTECH_NOT U256 ( .A(a[8]), .Z(n378) );
endmodule

