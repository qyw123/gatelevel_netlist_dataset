
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n85) );
  GTECH_XNOR2 U78 ( .A(n84), .B(n90), .Z(N154) );
  GTECH_XNOR2 U79 ( .A(n91), .B(n92), .Z(n90) );
  GTECH_NOT U80 ( .A(n86), .Z(n92) );
  GTECH_XNOR2 U81 ( .A(n93), .B(n88), .Z(n86) );
  GTECH_NOT U82 ( .A(n94), .Z(n88) );
  GTECH_NAND2 U83 ( .A(I_b[7]), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U84 ( .A(n89), .Z(n93) );
  GTECH_OAI22 U85 ( .A(n95), .B(n96), .C(n97), .D(n98), .Z(n89) );
  GTECH_AND2 U86 ( .A(n95), .B(n96), .Z(n97) );
  GTECH_NOT U87 ( .A(n99), .Z(n95) );
  GTECH_NOT U88 ( .A(n87), .Z(n91) );
  GTECH_OAI2N2 U89 ( .A(n100), .B(n101), .C(n102), .D(n103), .Z(n87) );
  GTECH_NAND2 U90 ( .A(n100), .B(n101), .Z(n103) );
  GTECH_NOT U91 ( .A(n104), .Z(n84) );
  GTECH_NAND2 U92 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_NOT U93 ( .A(n107), .Z(n105) );
  GTECH_XNOR2 U94 ( .A(n106), .B(n107), .Z(N153) );
  GTECH_XOR3 U95 ( .A(n108), .B(n100), .C(n102), .Z(n107) );
  GTECH_XOR3 U96 ( .A(n109), .B(n110), .C(n99), .Z(n102) );
  GTECH_OAI22 U97 ( .A(n111), .B(n112), .C(n113), .D(n114), .Z(n99) );
  GTECH_AND2 U98 ( .A(n111), .B(n112), .Z(n113) );
  GTECH_NOT U99 ( .A(n115), .Z(n111) );
  GTECH_NOT U100 ( .A(n98), .Z(n110) );
  GTECH_NAND2 U101 ( .A(I_b[7]), .B(I_a[6]), .Z(n98) );
  GTECH_NOT U102 ( .A(n96), .Z(n109) );
  GTECH_NAND2 U103 ( .A(I_a[7]), .B(I_b[6]), .Z(n96) );
  GTECH_ADD_ABC U104 ( .A(n116), .B(n117), .C(n118), .COUT(n100) );
  GTECH_NOT U105 ( .A(n119), .Z(n118) );
  GTECH_XNOR2 U106 ( .A(n120), .B(n121), .Z(n117) );
  GTECH_NAND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n121) );
  GTECH_NOT U108 ( .A(n101), .Z(n108) );
  GTECH_NAND2 U109 ( .A(I_a[7]), .B(n122), .Z(n101) );
  GTECH_NOT U110 ( .A(n123), .Z(n106) );
  GTECH_NAND2 U111 ( .A(n124), .B(n125), .Z(n123) );
  GTECH_NOT U112 ( .A(n126), .Z(n125) );
  GTECH_XNOR2 U113 ( .A(n126), .B(n124), .Z(N152) );
  GTECH_XOR4 U114 ( .A(n120), .B(n127), .C(n116), .D(n119), .Z(n124) );
  GTECH_XOR3 U115 ( .A(n128), .B(n129), .C(n115), .Z(n119) );
  GTECH_OAI22 U116 ( .A(n130), .B(n131), .C(n132), .D(n133), .Z(n115) );
  GTECH_AND2 U117 ( .A(n130), .B(n131), .Z(n132) );
  GTECH_NOT U118 ( .A(n134), .Z(n130) );
  GTECH_NOT U119 ( .A(n114), .Z(n129) );
  GTECH_NAND2 U120 ( .A(I_b[7]), .B(I_a[5]), .Z(n114) );
  GTECH_NOT U121 ( .A(n112), .Z(n128) );
  GTECH_NAND2 U122 ( .A(I_b[6]), .B(I_a[6]), .Z(n112) );
  GTECH_ADD_ABC U123 ( .A(n135), .B(n136), .C(n137), .COUT(n116) );
  GTECH_NOT U124 ( .A(n138), .Z(n137) );
  GTECH_XOR3 U125 ( .A(n139), .B(n140), .C(n141), .Z(n136) );
  GTECH_NOT U126 ( .A(n142), .Z(n139) );
  GTECH_AND2 U127 ( .A(I_a[7]), .B(I_b[5]), .Z(n127) );
  GTECH_NOT U128 ( .A(n122), .Z(n120) );
  GTECH_OAI22 U129 ( .A(n141), .B(n142), .C(n143), .D(n144), .Z(n122) );
  GTECH_AND2 U130 ( .A(n141), .B(n142), .Z(n143) );
  GTECH_NOT U131 ( .A(n145), .Z(n141) );
  GTECH_ADD_ABC U132 ( .A(n146), .B(n147), .C(n148), .COUT(n126) );
  GTECH_NOT U133 ( .A(n149), .Z(n148) );
  GTECH_OA22 U134 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n147) );
  GTECH_OA21 U135 ( .A(n154), .B(n155), .C(n156), .Z(n146) );
  GTECH_AO21 U136 ( .A(n154), .B(n155), .C(n157), .Z(n156) );
  GTECH_XOR3 U137 ( .A(n158), .B(n149), .C(n159), .Z(N151) );
  GTECH_OA21 U138 ( .A(n154), .B(n155), .C(n160), .Z(n159) );
  GTECH_AO21 U139 ( .A(n154), .B(n155), .C(n157), .Z(n160) );
  GTECH_XOR3 U140 ( .A(n138), .B(n135), .C(n161), .Z(n149) );
  GTECH_XOR3 U141 ( .A(n140), .B(n145), .C(n142), .Z(n161) );
  GTECH_NAND2 U142 ( .A(I_a[7]), .B(I_b[4]), .Z(n142) );
  GTECH_OAI22 U143 ( .A(n162), .B(n163), .C(n164), .D(n165), .Z(n145) );
  GTECH_AND2 U144 ( .A(n162), .B(n163), .Z(n164) );
  GTECH_NOT U145 ( .A(n144), .Z(n140) );
  GTECH_NAND2 U146 ( .A(I_a[6]), .B(I_b[5]), .Z(n144) );
  GTECH_ADD_ABC U147 ( .A(n166), .B(n167), .C(n168), .COUT(n135) );
  GTECH_NOT U148 ( .A(n169), .Z(n168) );
  GTECH_XOR3 U149 ( .A(n170), .B(n171), .C(n162), .Z(n167) );
  GTECH_NOT U150 ( .A(n172), .Z(n162) );
  GTECH_XOR3 U151 ( .A(n173), .B(n174), .C(n134), .Z(n138) );
  GTECH_OAI22 U152 ( .A(n175), .B(n176), .C(n177), .D(n178), .Z(n134) );
  GTECH_AND2 U153 ( .A(n175), .B(n176), .Z(n177) );
  GTECH_NOT U154 ( .A(n179), .Z(n175) );
  GTECH_NOT U155 ( .A(n133), .Z(n174) );
  GTECH_NAND2 U156 ( .A(I_b[7]), .B(I_a[4]), .Z(n133) );
  GTECH_NOT U157 ( .A(n131), .Z(n173) );
  GTECH_NAND2 U158 ( .A(I_b[6]), .B(I_a[5]), .Z(n131) );
  GTECH_OA22 U159 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n158) );
  GTECH_NOT U160 ( .A(I_a[7]), .Z(n151) );
  GTECH_XOR3 U161 ( .A(n154), .B(n180), .C(n157), .Z(N150) );
  GTECH_XOR3 U162 ( .A(n181), .B(n169), .C(n166), .Z(n157) );
  GTECH_ADD_ABC U163 ( .A(n182), .B(n183), .C(n184), .COUT(n166) );
  GTECH_NOT U164 ( .A(n185), .Z(n184) );
  GTECH_XOR3 U165 ( .A(n186), .B(n187), .C(n188), .Z(n183) );
  GTECH_XOR3 U166 ( .A(n189), .B(n190), .C(n179), .Z(n169) );
  GTECH_OAI22 U167 ( .A(n191), .B(n192), .C(n193), .D(n194), .Z(n179) );
  GTECH_AND2 U168 ( .A(n191), .B(n192), .Z(n193) );
  GTECH_NOT U169 ( .A(n195), .Z(n191) );
  GTECH_NOT U170 ( .A(n178), .Z(n190) );
  GTECH_NAND2 U171 ( .A(I_b[7]), .B(I_a[3]), .Z(n178) );
  GTECH_NOT U172 ( .A(n176), .Z(n189) );
  GTECH_NAND2 U173 ( .A(I_b[6]), .B(I_a[4]), .Z(n176) );
  GTECH_XOR3 U174 ( .A(n171), .B(n172), .C(n170), .Z(n181) );
  GTECH_NOT U175 ( .A(n163), .Z(n170) );
  GTECH_NAND2 U176 ( .A(I_a[6]), .B(I_b[4]), .Z(n163) );
  GTECH_OAI22 U177 ( .A(n188), .B(n196), .C(n197), .D(n198), .Z(n172) );
  GTECH_AND2 U178 ( .A(n188), .B(n196), .Z(n197) );
  GTECH_NOT U179 ( .A(n199), .Z(n188) );
  GTECH_NOT U180 ( .A(n165), .Z(n171) );
  GTECH_NAND2 U181 ( .A(I_a[5]), .B(I_b[5]), .Z(n165) );
  GTECH_NOT U182 ( .A(n155), .Z(n180) );
  GTECH_XNOR2 U183 ( .A(n152), .B(n153), .Z(n155) );
  GTECH_XNOR2 U184 ( .A(n150), .B(n200), .Z(n153) );
  GTECH_NAND2 U185 ( .A(I_a[7]), .B(I_b[3]), .Z(n200) );
  GTECH_OA21 U186 ( .A(n201), .B(n202), .C(n203), .Z(n150) );
  GTECH_AO21 U187 ( .A(n201), .B(n202), .C(n204), .Z(n203) );
  GTECH_NOT U188 ( .A(n205), .Z(n201) );
  GTECH_AOI2N2 U189 ( .A(n206), .B(n207), .C(n208), .D(n209), .Z(n152) );
  GTECH_NAND2 U190 ( .A(n208), .B(n209), .Z(n207) );
  GTECH_OA21 U191 ( .A(n210), .B(n211), .C(n212), .Z(n154) );
  GTECH_AO21 U192 ( .A(n210), .B(n211), .C(n213), .Z(n212) );
  GTECH_XOR3 U193 ( .A(n210), .B(n214), .C(n213), .Z(N149) );
  GTECH_XOR3 U194 ( .A(n215), .B(n185), .C(n182), .Z(n213) );
  GTECH_ADD_ABC U195 ( .A(n216), .B(n217), .C(n218), .COUT(n182) );
  GTECH_XOR3 U196 ( .A(n219), .B(n220), .C(n221), .Z(n217) );
  GTECH_OA21 U197 ( .A(n222), .B(n223), .C(n224), .Z(n216) );
  GTECH_AO21 U198 ( .A(n222), .B(n223), .C(n225), .Z(n224) );
  GTECH_XOR3 U199 ( .A(n226), .B(n227), .C(n195), .Z(n185) );
  GTECH_AO21 U200 ( .A(n228), .B(n229), .C(n230), .Z(n195) );
  GTECH_NOT U201 ( .A(n231), .Z(n230) );
  GTECH_NOT U202 ( .A(n194), .Z(n227) );
  GTECH_NAND2 U203 ( .A(I_b[7]), .B(I_a[2]), .Z(n194) );
  GTECH_NOT U204 ( .A(n192), .Z(n226) );
  GTECH_NAND2 U205 ( .A(I_b[6]), .B(I_a[3]), .Z(n192) );
  GTECH_XOR3 U206 ( .A(n187), .B(n199), .C(n186), .Z(n215) );
  GTECH_NOT U207 ( .A(n196), .Z(n186) );
  GTECH_NAND2 U208 ( .A(I_a[5]), .B(I_b[4]), .Z(n196) );
  GTECH_OAI22 U209 ( .A(n221), .B(n232), .C(n233), .D(n234), .Z(n199) );
  GTECH_AND2 U210 ( .A(n221), .B(n232), .Z(n233) );
  GTECH_NOT U211 ( .A(n235), .Z(n221) );
  GTECH_NOT U212 ( .A(n198), .Z(n187) );
  GTECH_NAND2 U213 ( .A(I_b[5]), .B(I_a[4]), .Z(n198) );
  GTECH_NOT U214 ( .A(n211), .Z(n214) );
  GTECH_XOR3 U215 ( .A(n236), .B(n208), .C(n206), .Z(n211) );
  GTECH_XOR3 U216 ( .A(n237), .B(n238), .C(n205), .Z(n206) );
  GTECH_OAI22 U217 ( .A(n239), .B(n240), .C(n241), .D(n242), .Z(n205) );
  GTECH_AND2 U218 ( .A(n239), .B(n240), .Z(n241) );
  GTECH_NOT U219 ( .A(n243), .Z(n239) );
  GTECH_NOT U220 ( .A(n204), .Z(n238) );
  GTECH_NAND2 U221 ( .A(I_a[6]), .B(I_b[3]), .Z(n204) );
  GTECH_NOT U222 ( .A(n202), .Z(n237) );
  GTECH_NAND2 U223 ( .A(I_a[7]), .B(I_b[2]), .Z(n202) );
  GTECH_ADD_ABC U224 ( .A(n244), .B(n245), .C(n246), .COUT(n208) );
  GTECH_XNOR2 U225 ( .A(n247), .B(n248), .Z(n245) );
  GTECH_NAND2 U226 ( .A(I_a[7]), .B(I_b[1]), .Z(n248) );
  GTECH_NOT U227 ( .A(n209), .Z(n236) );
  GTECH_NAND2 U228 ( .A(I_a[7]), .B(n249), .Z(n209) );
  GTECH_ADD_ABC U229 ( .A(n250), .B(n251), .C(n252), .COUT(n210) );
  GTECH_XOR3 U230 ( .A(n244), .B(n253), .C(n246), .Z(n251) );
  GTECH_NOT U231 ( .A(n254), .Z(n246) );
  GTECH_XOR3 U232 ( .A(n255), .B(n252), .C(n250), .Z(N148) );
  GTECH_ADD_ABC U233 ( .A(n256), .B(n257), .C(n258), .COUT(n250) );
  GTECH_NOT U234 ( .A(n259), .Z(n258) );
  GTECH_XOR3 U235 ( .A(n260), .B(n261), .C(n262), .Z(n257) );
  GTECH_NOT U236 ( .A(n263), .Z(n261) );
  GTECH_XOR3 U237 ( .A(n264), .B(n218), .C(n265), .Z(n252) );
  GTECH_OAI22 U238 ( .A(n222), .B(n223), .C(n266), .D(n225), .Z(n265) );
  GTECH_AND2 U239 ( .A(n222), .B(n223), .Z(n266) );
  GTECH_XOR3 U240 ( .A(n229), .B(n228), .C(n231), .Z(n218) );
  GTECH_NAND3 U241 ( .A(I_b[6]), .B(I_a[1]), .C(n267), .Z(n231) );
  GTECH_NOT U242 ( .A(n268), .Z(n228) );
  GTECH_NAND2 U243 ( .A(I_b[7]), .B(I_a[1]), .Z(n268) );
  GTECH_NOT U244 ( .A(n269), .Z(n229) );
  GTECH_NAND2 U245 ( .A(I_b[6]), .B(I_a[2]), .Z(n269) );
  GTECH_XOR3 U246 ( .A(n220), .B(n235), .C(n219), .Z(n264) );
  GTECH_NOT U247 ( .A(n232), .Z(n219) );
  GTECH_NAND2 U248 ( .A(I_b[4]), .B(I_a[4]), .Z(n232) );
  GTECH_OAI22 U249 ( .A(n270), .B(n271), .C(n272), .D(n273), .Z(n235) );
  GTECH_AND2 U250 ( .A(n270), .B(n271), .Z(n272) );
  GTECH_NOT U251 ( .A(n274), .Z(n270) );
  GTECH_NOT U252 ( .A(n234), .Z(n220) );
  GTECH_NAND2 U253 ( .A(I_b[5]), .B(I_a[3]), .Z(n234) );
  GTECH_XOR3 U254 ( .A(n253), .B(n254), .C(n244), .Z(n255) );
  GTECH_ADD_ABC U255 ( .A(n260), .B(n275), .C(n262), .COUT(n244) );
  GTECH_NOT U256 ( .A(n276), .Z(n262) );
  GTECH_XOR3 U257 ( .A(n277), .B(n278), .C(n279), .Z(n275) );
  GTECH_XOR3 U258 ( .A(n280), .B(n281), .C(n243), .Z(n254) );
  GTECH_OAI22 U259 ( .A(n282), .B(n283), .C(n284), .D(n285), .Z(n243) );
  GTECH_AND2 U260 ( .A(n282), .B(n283), .Z(n284) );
  GTECH_NOT U261 ( .A(n286), .Z(n282) );
  GTECH_NOT U262 ( .A(n242), .Z(n281) );
  GTECH_NAND2 U263 ( .A(I_a[5]), .B(I_b[3]), .Z(n242) );
  GTECH_NOT U264 ( .A(n240), .Z(n280) );
  GTECH_NAND2 U265 ( .A(I_a[6]), .B(I_b[2]), .Z(n240) );
  GTECH_XNOR2 U266 ( .A(n247), .B(n287), .Z(n253) );
  GTECH_NAND2 U267 ( .A(I_a[7]), .B(I_b[1]), .Z(n287) );
  GTECH_NOT U268 ( .A(n249), .Z(n247) );
  GTECH_OAI22 U269 ( .A(n279), .B(n288), .C(n289), .D(n290), .Z(n249) );
  GTECH_AND2 U270 ( .A(n279), .B(n288), .Z(n289) );
  GTECH_NOT U271 ( .A(n291), .Z(n279) );
  GTECH_XOR3 U272 ( .A(n259), .B(n256), .C(n292), .Z(N147) );
  GTECH_XOR3 U273 ( .A(n276), .B(n260), .C(n263), .Z(n292) );
  GTECH_XOR3 U274 ( .A(n277), .B(n278), .C(n291), .Z(n263) );
  GTECH_OAI22 U275 ( .A(n293), .B(n294), .C(n295), .D(n296), .Z(n291) );
  GTECH_AND2 U276 ( .A(n293), .B(n294), .Z(n295) );
  GTECH_NOT U277 ( .A(n290), .Z(n278) );
  GTECH_NAND2 U278 ( .A(I_a[6]), .B(I_b[1]), .Z(n290) );
  GTECH_NOT U279 ( .A(n288), .Z(n277) );
  GTECH_NAND2 U280 ( .A(I_a[7]), .B(I_b[0]), .Z(n288) );
  GTECH_ADD_ABC U281 ( .A(n297), .B(n298), .C(n299), .COUT(n260) );
  GTECH_XOR3 U282 ( .A(n300), .B(n301), .C(n293), .Z(n298) );
  GTECH_NOT U283 ( .A(n302), .Z(n293) );
  GTECH_XOR3 U284 ( .A(n303), .B(n304), .C(n286), .Z(n276) );
  GTECH_OAI22 U285 ( .A(n305), .B(n306), .C(n307), .D(n308), .Z(n286) );
  GTECH_AND2 U286 ( .A(n305), .B(n306), .Z(n307) );
  GTECH_NOT U287 ( .A(n309), .Z(n305) );
  GTECH_NOT U288 ( .A(n285), .Z(n304) );
  GTECH_NAND2 U289 ( .A(I_b[3]), .B(I_a[4]), .Z(n285) );
  GTECH_NOT U290 ( .A(n283), .Z(n303) );
  GTECH_NAND2 U291 ( .A(I_a[5]), .B(I_b[2]), .Z(n283) );
  GTECH_ADD_ABC U292 ( .A(n310), .B(n311), .C(n312), .COUT(n256) );
  GTECH_XOR3 U293 ( .A(n297), .B(n313), .C(n299), .Z(n311) );
  GTECH_NOT U294 ( .A(n314), .Z(n299) );
  GTECH_OA21 U295 ( .A(n315), .B(n316), .C(n317), .Z(n310) );
  GTECH_AO21 U296 ( .A(n315), .B(n316), .C(n318), .Z(n317) );
  GTECH_XOR3 U297 ( .A(n319), .B(n223), .C(n222), .Z(n259) );
  GTECH_XNOR2 U298 ( .A(n267), .B(n320), .Z(n222) );
  GTECH_AND2 U299 ( .A(I_b[6]), .B(I_a[1]), .Z(n320) );
  GTECH_NOT U300 ( .A(n321), .Z(n267) );
  GTECH_NAND2 U301 ( .A(I_b[7]), .B(I_a[0]), .Z(n321) );
  GTECH_NOT U302 ( .A(n322), .Z(n223) );
  GTECH_XOR3 U303 ( .A(n323), .B(n324), .C(n274), .Z(n322) );
  GTECH_AO21 U304 ( .A(n325), .B(n326), .C(n327), .Z(n274) );
  GTECH_NOT U305 ( .A(n328), .Z(n327) );
  GTECH_NOT U306 ( .A(n273), .Z(n324) );
  GTECH_NAND2 U307 ( .A(I_b[5]), .B(I_a[2]), .Z(n273) );
  GTECH_NOT U308 ( .A(n271), .Z(n323) );
  GTECH_NAND2 U309 ( .A(I_b[4]), .B(I_a[3]), .Z(n271) );
  GTECH_NOT U310 ( .A(n225), .Z(n319) );
  GTECH_NAND3 U311 ( .A(I_a[0]), .B(n329), .C(I_b[6]), .Z(n225) );
  GTECH_XOR3 U312 ( .A(n330), .B(n312), .C(n331), .Z(N146) );
  GTECH_OA21 U313 ( .A(n315), .B(n316), .C(n332), .Z(n331) );
  GTECH_AO21 U314 ( .A(n315), .B(n316), .C(n318), .Z(n332) );
  GTECH_XNOR2 U315 ( .A(n333), .B(n329), .Z(n312) );
  GTECH_NOT U316 ( .A(n334), .Z(n329) );
  GTECH_XOR3 U317 ( .A(n326), .B(n325), .C(n328), .Z(n334) );
  GTECH_NAND3 U318 ( .A(I_b[4]), .B(I_a[1]), .C(n335), .Z(n328) );
  GTECH_NOT U319 ( .A(n336), .Z(n325) );
  GTECH_NAND2 U320 ( .A(I_b[5]), .B(I_a[1]), .Z(n336) );
  GTECH_NOT U321 ( .A(n337), .Z(n326) );
  GTECH_NAND2 U322 ( .A(I_b[4]), .B(I_a[2]), .Z(n337) );
  GTECH_AND2 U323 ( .A(I_b[6]), .B(I_a[0]), .Z(n333) );
  GTECH_XOR3 U324 ( .A(n313), .B(n314), .C(n297), .Z(n330) );
  GTECH_ADD_ABC U325 ( .A(n338), .B(n339), .C(n340), .COUT(n297) );
  GTECH_NOT U326 ( .A(n341), .Z(n340) );
  GTECH_XOR3 U327 ( .A(n342), .B(n343), .C(n344), .Z(n339) );
  GTECH_XOR3 U328 ( .A(n345), .B(n346), .C(n309), .Z(n314) );
  GTECH_OAI22 U329 ( .A(n347), .B(n348), .C(n349), .D(n350), .Z(n309) );
  GTECH_AND2 U330 ( .A(n347), .B(n348), .Z(n349) );
  GTECH_NOT U331 ( .A(n351), .Z(n347) );
  GTECH_NOT U332 ( .A(n308), .Z(n346) );
  GTECH_NAND2 U333 ( .A(I_b[3]), .B(I_a[3]), .Z(n308) );
  GTECH_NOT U334 ( .A(n306), .Z(n345) );
  GTECH_NAND2 U335 ( .A(I_b[2]), .B(I_a[4]), .Z(n306) );
  GTECH_NOT U336 ( .A(n352), .Z(n313) );
  GTECH_XOR3 U337 ( .A(n300), .B(n301), .C(n302), .Z(n352) );
  GTECH_OAI22 U338 ( .A(n344), .B(n353), .C(n354), .D(n355), .Z(n302) );
  GTECH_AND2 U339 ( .A(n344), .B(n353), .Z(n354) );
  GTECH_NOT U340 ( .A(n356), .Z(n344) );
  GTECH_NOT U341 ( .A(n296), .Z(n301) );
  GTECH_NAND2 U342 ( .A(I_a[5]), .B(I_b[1]), .Z(n296) );
  GTECH_NOT U343 ( .A(n294), .Z(n300) );
  GTECH_NAND2 U344 ( .A(I_a[6]), .B(I_b[0]), .Z(n294) );
  GTECH_XOR3 U345 ( .A(n357), .B(n316), .C(n315), .Z(N145) );
  GTECH_XNOR2 U346 ( .A(n335), .B(n358), .Z(n315) );
  GTECH_AND2 U347 ( .A(I_b[4]), .B(I_a[1]), .Z(n358) );
  GTECH_NOT U348 ( .A(n359), .Z(n335) );
  GTECH_NAND2 U349 ( .A(I_b[5]), .B(I_a[0]), .Z(n359) );
  GTECH_XOR3 U350 ( .A(n360), .B(n341), .C(n338), .Z(n316) );
  GTECH_ADD_ABC U351 ( .A(n361), .B(n362), .C(n363), .COUT(n338) );
  GTECH_XOR3 U352 ( .A(n364), .B(n365), .C(n366), .Z(n362) );
  GTECH_OA21 U353 ( .A(n367), .B(n368), .C(n369), .Z(n361) );
  GTECH_AO21 U354 ( .A(n367), .B(n368), .C(n370), .Z(n369) );
  GTECH_XOR3 U355 ( .A(n371), .B(n372), .C(n351), .Z(n341) );
  GTECH_AO21 U356 ( .A(n373), .B(n374), .C(n375), .Z(n351) );
  GTECH_NOT U357 ( .A(n376), .Z(n375) );
  GTECH_NOT U358 ( .A(n350), .Z(n372) );
  GTECH_NAND2 U359 ( .A(I_b[3]), .B(I_a[2]), .Z(n350) );
  GTECH_NOT U360 ( .A(n348), .Z(n371) );
  GTECH_NAND2 U361 ( .A(I_b[2]), .B(I_a[3]), .Z(n348) );
  GTECH_XOR3 U362 ( .A(n343), .B(n356), .C(n342), .Z(n360) );
  GTECH_NOT U363 ( .A(n353), .Z(n342) );
  GTECH_NAND2 U364 ( .A(I_a[5]), .B(I_b[0]), .Z(n353) );
  GTECH_OAI22 U365 ( .A(n366), .B(n377), .C(n378), .D(n379), .Z(n356) );
  GTECH_AND2 U366 ( .A(n366), .B(n377), .Z(n378) );
  GTECH_NOT U367 ( .A(n380), .Z(n366) );
  GTECH_NOT U368 ( .A(n355), .Z(n343) );
  GTECH_NAND2 U369 ( .A(I_a[4]), .B(I_b[1]), .Z(n355) );
  GTECH_NOT U370 ( .A(n318), .Z(n357) );
  GTECH_NAND3 U371 ( .A(I_a[0]), .B(n381), .C(I_b[4]), .Z(n318) );
  GTECH_NOT U372 ( .A(n382), .Z(n381) );
  GTECH_XNOR2 U373 ( .A(n383), .B(n382), .Z(N144) );
  GTECH_XOR3 U374 ( .A(n384), .B(n363), .C(n385), .Z(n382) );
  GTECH_OAI22 U375 ( .A(n367), .B(n368), .C(n386), .D(n370), .Z(n385) );
  GTECH_AND2 U376 ( .A(n367), .B(n368), .Z(n386) );
  GTECH_XOR3 U377 ( .A(n374), .B(n373), .C(n376), .Z(n363) );
  GTECH_NAND3 U378 ( .A(I_b[2]), .B(I_a[1]), .C(n387), .Z(n376) );
  GTECH_NOT U379 ( .A(n388), .Z(n373) );
  GTECH_NAND2 U380 ( .A(I_b[3]), .B(I_a[1]), .Z(n388) );
  GTECH_NOT U381 ( .A(n389), .Z(n374) );
  GTECH_NAND2 U382 ( .A(I_b[2]), .B(I_a[2]), .Z(n389) );
  GTECH_XOR3 U383 ( .A(n365), .B(n380), .C(n364), .Z(n384) );
  GTECH_NOT U384 ( .A(n377), .Z(n364) );
  GTECH_NAND2 U385 ( .A(I_a[4]), .B(I_b[0]), .Z(n377) );
  GTECH_OAI22 U386 ( .A(n390), .B(n391), .C(n392), .D(n393), .Z(n380) );
  GTECH_AND2 U387 ( .A(n390), .B(n391), .Z(n392) );
  GTECH_NOT U388 ( .A(n394), .Z(n390) );
  GTECH_NOT U389 ( .A(n379), .Z(n365) );
  GTECH_NAND2 U390 ( .A(I_a[3]), .B(I_b[1]), .Z(n379) );
  GTECH_AND2 U391 ( .A(I_b[4]), .B(I_a[0]), .Z(n383) );
  GTECH_XOR3 U392 ( .A(n395), .B(n368), .C(n367), .Z(N143) );
  GTECH_XNOR2 U393 ( .A(n387), .B(n396), .Z(n367) );
  GTECH_AND2 U394 ( .A(I_b[2]), .B(I_a[1]), .Z(n396) );
  GTECH_NOT U395 ( .A(n397), .Z(n387) );
  GTECH_NAND2 U396 ( .A(I_b[3]), .B(I_a[0]), .Z(n397) );
  GTECH_NOT U397 ( .A(n398), .Z(n368) );
  GTECH_XOR3 U398 ( .A(n399), .B(n400), .C(n394), .Z(n398) );
  GTECH_AO21 U399 ( .A(n401), .B(n402), .C(n403), .Z(n394) );
  GTECH_NOT U400 ( .A(n404), .Z(n403) );
  GTECH_NOT U401 ( .A(n393), .Z(n400) );
  GTECH_NAND2 U402 ( .A(I_b[1]), .B(I_a[2]), .Z(n393) );
  GTECH_NOT U403 ( .A(n391), .Z(n399) );
  GTECH_NAND2 U404 ( .A(I_b[0]), .B(I_a[3]), .Z(n391) );
  GTECH_NOT U405 ( .A(n370), .Z(n395) );
  GTECH_NAND3 U406 ( .A(I_a[0]), .B(n405), .C(I_b[2]), .Z(n370) );
  GTECH_NOT U407 ( .A(n406), .Z(n405) );
  GTECH_XNOR2 U408 ( .A(n407), .B(n406), .Z(N142) );
  GTECH_XOR3 U409 ( .A(n401), .B(n402), .C(n404), .Z(n406) );
  GTECH_NAND3 U410 ( .A(n408), .B(I_b[0]), .C(I_a[1]), .Z(n404) );
  GTECH_NOT U411 ( .A(n409), .Z(n402) );
  GTECH_NAND2 U412 ( .A(I_a[1]), .B(I_b[1]), .Z(n409) );
  GTECH_NOT U413 ( .A(n410), .Z(n401) );
  GTECH_NAND2 U414 ( .A(I_b[0]), .B(I_a[2]), .Z(n410) );
  GTECH_AND2 U415 ( .A(I_b[2]), .B(I_a[0]), .Z(n407) );
  GTECH_XNOR2 U416 ( .A(n408), .B(n411), .Z(N141) );
  GTECH_NAND2 U417 ( .A(I_a[1]), .B(I_b[0]), .Z(n411) );
  GTECH_NOT U418 ( .A(n412), .Z(n408) );
  GTECH_NAND2 U419 ( .A(I_a[0]), .B(I_b[1]), .Z(n412) );
  GTECH_AND2 U420 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

