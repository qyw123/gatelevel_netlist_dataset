
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI21 U82 ( .A(n93), .B(n94), .C(n95), .Z(n87) );
  GTECH_OAI21 U83 ( .A(n96), .B(n97), .C(n98), .Z(n95) );
  GTECH_NOT U84 ( .A(n93), .Z(n97) );
  GTECH_XOR2 U85 ( .A(n90), .B(n99), .Z(n86) );
  GTECH_NOT U86 ( .A(n89), .Z(n99) );
  GTECH_OAI21 U87 ( .A(n100), .B(n101), .C(n102), .Z(n89) );
  GTECH_OAI21 U88 ( .A(n103), .B(n104), .C(n105), .Z(n102) );
  GTECH_NOT U89 ( .A(n104), .Z(n100) );
  GTECH_NAND2 U90 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U91 ( .A(n106), .Z(n84) );
  GTECH_NAND2 U92 ( .A(n107), .B(n108), .Z(n106) );
  GTECH_XOR2 U93 ( .A(n108), .B(n107), .Z(N153) );
  GTECH_NOT U94 ( .A(n109), .Z(n107) );
  GTECH_XOR3 U95 ( .A(n96), .B(n93), .C(n98), .Z(n109) );
  GTECH_XOR3 U96 ( .A(n103), .B(n105), .C(n104), .Z(n98) );
  GTECH_OAI21 U97 ( .A(n110), .B(n111), .C(n112), .Z(n104) );
  GTECH_OAI21 U98 ( .A(n113), .B(n114), .C(n115), .Z(n112) );
  GTECH_NOT U99 ( .A(n114), .Z(n110) );
  GTECH_NOT U100 ( .A(n116), .Z(n105) );
  GTECH_NAND2 U101 ( .A(I_b[7]), .B(I_a[6]), .Z(n116) );
  GTECH_NOT U102 ( .A(n101), .Z(n103) );
  GTECH_NAND2 U103 ( .A(I_a[7]), .B(I_b[6]), .Z(n101) );
  GTECH_ADD_ABC U104 ( .A(n117), .B(n118), .C(n119), .COUT(n93) );
  GTECH_NOT U105 ( .A(n120), .Z(n119) );
  GTECH_XOR2 U106 ( .A(n121), .B(n122), .Z(n118) );
  GTECH_AND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n122) );
  GTECH_NOT U108 ( .A(n123), .Z(n121) );
  GTECH_NOT U109 ( .A(n94), .Z(n96) );
  GTECH_NAND2 U110 ( .A(I_a[7]), .B(n123), .Z(n94) );
  GTECH_NOT U111 ( .A(n124), .Z(n108) );
  GTECH_NAND2 U112 ( .A(n125), .B(n126), .Z(n124) );
  GTECH_NOT U113 ( .A(n127), .Z(n126) );
  GTECH_XOR2 U114 ( .A(n127), .B(n128), .Z(N152) );
  GTECH_NOT U115 ( .A(n125), .Z(n128) );
  GTECH_XNOR4 U116 ( .A(n129), .B(n120), .C(n123), .D(n117), .Z(n125) );
  GTECH_ADD_ABC U117 ( .A(n130), .B(n131), .C(n132), .COUT(n117) );
  GTECH_NOT U118 ( .A(n133), .Z(n132) );
  GTECH_XOR3 U119 ( .A(n134), .B(n135), .C(n136), .Z(n131) );
  GTECH_OAI21 U120 ( .A(n136), .B(n137), .C(n138), .Z(n123) );
  GTECH_OAI21 U121 ( .A(n134), .B(n139), .C(n135), .Z(n138) );
  GTECH_NOT U122 ( .A(n139), .Z(n136) );
  GTECH_XOR3 U123 ( .A(n113), .B(n115), .C(n114), .Z(n120) );
  GTECH_OAI21 U124 ( .A(n140), .B(n141), .C(n142), .Z(n114) );
  GTECH_OAI21 U125 ( .A(n143), .B(n144), .C(n145), .Z(n142) );
  GTECH_NOT U126 ( .A(n144), .Z(n140) );
  GTECH_NOT U127 ( .A(n146), .Z(n115) );
  GTECH_NAND2 U128 ( .A(I_b[7]), .B(I_a[5]), .Z(n146) );
  GTECH_NOT U129 ( .A(n111), .Z(n113) );
  GTECH_NAND2 U130 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_AND2 U131 ( .A(I_a[7]), .B(I_b[5]), .Z(n129) );
  GTECH_ADD_ABC U132 ( .A(n147), .B(n148), .C(n149), .COUT(n127) );
  GTECH_NOT U133 ( .A(n150), .Z(n149) );
  GTECH_OA22 U134 ( .A(n151), .B(n152), .C(n153), .D(n154), .Z(n148) );
  GTECH_OA21 U135 ( .A(n155), .B(n156), .C(n157), .Z(n147) );
  GTECH_XOR3 U136 ( .A(n158), .B(n150), .C(n159), .Z(N151) );
  GTECH_OA21 U137 ( .A(n155), .B(n156), .C(n157), .Z(n159) );
  GTECH_OAI21 U138 ( .A(n160), .B(n161), .C(n162), .Z(n157) );
  GTECH_XOR2 U139 ( .A(n163), .B(n130), .Z(n150) );
  GTECH_ADD_ABC U140 ( .A(n164), .B(n165), .C(n166), .COUT(n130) );
  GTECH_NOT U141 ( .A(n167), .Z(n166) );
  GTECH_XOR3 U142 ( .A(n168), .B(n169), .C(n170), .Z(n165) );
  GTECH_XNOR4 U143 ( .A(n135), .B(n139), .C(n133), .D(n134), .Z(n163) );
  GTECH_NOT U144 ( .A(n137), .Z(n134) );
  GTECH_NAND2 U145 ( .A(I_a[7]), .B(I_b[4]), .Z(n137) );
  GTECH_XOR3 U146 ( .A(n143), .B(n145), .C(n144), .Z(n133) );
  GTECH_OAI21 U147 ( .A(n171), .B(n172), .C(n173), .Z(n144) );
  GTECH_OAI21 U148 ( .A(n174), .B(n175), .C(n176), .Z(n173) );
  GTECH_NOT U149 ( .A(n175), .Z(n171) );
  GTECH_NOT U150 ( .A(n177), .Z(n145) );
  GTECH_NAND2 U151 ( .A(I_b[7]), .B(I_a[4]), .Z(n177) );
  GTECH_NOT U152 ( .A(n141), .Z(n143) );
  GTECH_NAND2 U153 ( .A(I_b[6]), .B(I_a[5]), .Z(n141) );
  GTECH_OAI21 U154 ( .A(n170), .B(n178), .C(n179), .Z(n139) );
  GTECH_OAI21 U155 ( .A(n168), .B(n180), .C(n169), .Z(n179) );
  GTECH_NOT U156 ( .A(n180), .Z(n170) );
  GTECH_NOT U157 ( .A(n181), .Z(n135) );
  GTECH_NAND2 U158 ( .A(I_a[6]), .B(I_b[5]), .Z(n181) );
  GTECH_OA22 U159 ( .A(n151), .B(n152), .C(n153), .D(n154), .Z(n158) );
  GTECH_NOT U160 ( .A(n182), .Z(n154) );
  GTECH_NOT U161 ( .A(I_a[7]), .Z(n152) );
  GTECH_XOR3 U162 ( .A(n155), .B(n160), .C(n183), .Z(N150) );
  GTECH_NOT U163 ( .A(n162), .Z(n183) );
  GTECH_XOR2 U164 ( .A(n184), .B(n164), .Z(n162) );
  GTECH_ADD_ABC U165 ( .A(n185), .B(n186), .C(n187), .COUT(n164) );
  GTECH_NOT U166 ( .A(n188), .Z(n187) );
  GTECH_XOR3 U167 ( .A(n189), .B(n190), .C(n191), .Z(n186) );
  GTECH_XNOR4 U168 ( .A(n169), .B(n180), .C(n167), .D(n168), .Z(n184) );
  GTECH_NOT U169 ( .A(n178), .Z(n168) );
  GTECH_NAND2 U170 ( .A(I_a[6]), .B(I_b[4]), .Z(n178) );
  GTECH_XOR3 U171 ( .A(n174), .B(n176), .C(n175), .Z(n167) );
  GTECH_OAI21 U172 ( .A(n192), .B(n193), .C(n194), .Z(n175) );
  GTECH_OAI21 U173 ( .A(n195), .B(n196), .C(n197), .Z(n194) );
  GTECH_NOT U174 ( .A(n196), .Z(n192) );
  GTECH_NOT U175 ( .A(n198), .Z(n176) );
  GTECH_NAND2 U176 ( .A(I_b[7]), .B(I_a[3]), .Z(n198) );
  GTECH_NOT U177 ( .A(n172), .Z(n174) );
  GTECH_NAND2 U178 ( .A(I_b[6]), .B(I_a[4]), .Z(n172) );
  GTECH_OAI21 U179 ( .A(n191), .B(n199), .C(n200), .Z(n180) );
  GTECH_OAI21 U180 ( .A(n189), .B(n201), .C(n190), .Z(n200) );
  GTECH_NOT U181 ( .A(n201), .Z(n191) );
  GTECH_NOT U182 ( .A(n202), .Z(n169) );
  GTECH_NAND2 U183 ( .A(I_a[5]), .B(I_b[5]), .Z(n202) );
  GTECH_NOT U184 ( .A(n156), .Z(n160) );
  GTECH_XOR2 U185 ( .A(n182), .B(n153), .Z(n156) );
  GTECH_AOI2N2 U186 ( .A(n203), .B(n204), .C(n205), .D(n206), .Z(n153) );
  GTECH_NAND2 U187 ( .A(n205), .B(n206), .Z(n204) );
  GTECH_XOR2 U188 ( .A(n207), .B(n151), .Z(n182) );
  GTECH_AND2 U189 ( .A(n208), .B(n209), .Z(n151) );
  GTECH_OR_NOT U190 ( .A(n210), .B(n211), .Z(n209) );
  GTECH_OAI21 U191 ( .A(n212), .B(n211), .C(n213), .Z(n208) );
  GTECH_NAND2 U192 ( .A(I_a[7]), .B(I_b[3]), .Z(n207) );
  GTECH_NOT U193 ( .A(n161), .Z(n155) );
  GTECH_OAI21 U194 ( .A(n214), .B(n215), .C(n216), .Z(n161) );
  GTECH_OAI21 U195 ( .A(n217), .B(n218), .C(n219), .Z(n216) );
  GTECH_NOT U196 ( .A(n214), .Z(n218) );
  GTECH_XOR3 U197 ( .A(n214), .B(n217), .C(n220), .Z(N149) );
  GTECH_NOT U198 ( .A(n219), .Z(n220) );
  GTECH_XOR2 U199 ( .A(n221), .B(n185), .Z(n219) );
  GTECH_ADD_ABC U200 ( .A(n222), .B(n223), .C(n224), .COUT(n185) );
  GTECH_XOR3 U201 ( .A(n225), .B(n226), .C(n227), .Z(n223) );
  GTECH_OA21 U202 ( .A(n228), .B(n229), .C(n230), .Z(n222) );
  GTECH_XNOR4 U203 ( .A(n190), .B(n201), .C(n188), .D(n189), .Z(n221) );
  GTECH_NOT U204 ( .A(n199), .Z(n189) );
  GTECH_NAND2 U205 ( .A(I_a[5]), .B(I_b[4]), .Z(n199) );
  GTECH_XOR3 U206 ( .A(n195), .B(n197), .C(n196), .Z(n188) );
  GTECH_OAI21 U207 ( .A(n231), .B(n232), .C(n233), .Z(n196) );
  GTECH_NOT U208 ( .A(n234), .Z(n197) );
  GTECH_NAND2 U209 ( .A(I_b[7]), .B(I_a[2]), .Z(n234) );
  GTECH_NOT U210 ( .A(n193), .Z(n195) );
  GTECH_NAND2 U211 ( .A(I_b[6]), .B(I_a[3]), .Z(n193) );
  GTECH_OAI21 U212 ( .A(n227), .B(n235), .C(n236), .Z(n201) );
  GTECH_OAI21 U213 ( .A(n225), .B(n237), .C(n226), .Z(n236) );
  GTECH_NOT U214 ( .A(n237), .Z(n227) );
  GTECH_NOT U215 ( .A(n238), .Z(n190) );
  GTECH_NAND2 U216 ( .A(I_b[5]), .B(I_a[4]), .Z(n238) );
  GTECH_NOT U217 ( .A(n215), .Z(n217) );
  GTECH_XOR3 U218 ( .A(n239), .B(n205), .C(n203), .Z(n215) );
  GTECH_XOR3 U219 ( .A(n212), .B(n213), .C(n211), .Z(n203) );
  GTECH_OAI21 U220 ( .A(n240), .B(n241), .C(n242), .Z(n211) );
  GTECH_OAI21 U221 ( .A(n243), .B(n244), .C(n245), .Z(n242) );
  GTECH_NOT U222 ( .A(n244), .Z(n240) );
  GTECH_NOT U223 ( .A(n246), .Z(n213) );
  GTECH_NAND2 U224 ( .A(I_a[6]), .B(I_b[3]), .Z(n246) );
  GTECH_NOT U225 ( .A(n210), .Z(n212) );
  GTECH_NAND2 U226 ( .A(I_a[7]), .B(I_b[2]), .Z(n210) );
  GTECH_ADD_ABC U227 ( .A(n247), .B(n248), .C(n249), .COUT(n205) );
  GTECH_XOR2 U228 ( .A(n250), .B(n251), .Z(n248) );
  GTECH_AND2 U229 ( .A(I_a[7]), .B(I_b[1]), .Z(n251) );
  GTECH_NOT U230 ( .A(n206), .Z(n239) );
  GTECH_NAND2 U231 ( .A(I_a[7]), .B(n252), .Z(n206) );
  GTECH_ADD_ABC U232 ( .A(n253), .B(n254), .C(n255), .COUT(n214) );
  GTECH_XOR3 U233 ( .A(n247), .B(n256), .C(n249), .Z(n254) );
  GTECH_NOT U234 ( .A(n257), .Z(n249) );
  GTECH_XOR3 U235 ( .A(n258), .B(n255), .C(n253), .Z(N148) );
  GTECH_ADD_ABC U236 ( .A(n259), .B(n260), .C(n261), .COUT(n253) );
  GTECH_NOT U237 ( .A(n262), .Z(n261) );
  GTECH_XOR3 U238 ( .A(n263), .B(n264), .C(n265), .Z(n260) );
  GTECH_XOR2 U239 ( .A(n266), .B(n267), .Z(n255) );
  GTECH_OA21 U240 ( .A(n228), .B(n229), .C(n230), .Z(n267) );
  GTECH_OAI21 U241 ( .A(n268), .B(n269), .C(n270), .Z(n230) );
  GTECH_NOT U242 ( .A(n228), .Z(n269) );
  GTECH_XNOR4 U243 ( .A(n226), .B(n237), .C(n224), .D(n225), .Z(n266) );
  GTECH_NOT U244 ( .A(n235), .Z(n225) );
  GTECH_NAND2 U245 ( .A(I_b[4]), .B(I_a[4]), .Z(n235) );
  GTECH_XOR3 U246 ( .A(n271), .B(n272), .C(n233), .Z(n224) );
  GTECH_NAND3 U247 ( .A(I_b[6]), .B(I_a[1]), .C(n273), .Z(n233) );
  GTECH_NOT U248 ( .A(n232), .Z(n272) );
  GTECH_NAND2 U249 ( .A(I_b[7]), .B(I_a[1]), .Z(n232) );
  GTECH_NOT U250 ( .A(n231), .Z(n271) );
  GTECH_NAND2 U251 ( .A(I_b[6]), .B(I_a[2]), .Z(n231) );
  GTECH_OAI21 U252 ( .A(n274), .B(n275), .C(n276), .Z(n237) );
  GTECH_OAI21 U253 ( .A(n277), .B(n278), .C(n279), .Z(n276) );
  GTECH_NOT U254 ( .A(n278), .Z(n274) );
  GTECH_NOT U255 ( .A(n280), .Z(n226) );
  GTECH_NAND2 U256 ( .A(I_b[5]), .B(I_a[3]), .Z(n280) );
  GTECH_XOR3 U257 ( .A(n256), .B(n257), .C(n247), .Z(n258) );
  GTECH_ADD_ABC U258 ( .A(n263), .B(n281), .C(n265), .COUT(n247) );
  GTECH_NOT U259 ( .A(n282), .Z(n265) );
  GTECH_XOR3 U260 ( .A(n283), .B(n284), .C(n285), .Z(n281) );
  GTECH_XOR3 U261 ( .A(n243), .B(n245), .C(n244), .Z(n257) );
  GTECH_OAI21 U262 ( .A(n286), .B(n287), .C(n288), .Z(n244) );
  GTECH_OAI21 U263 ( .A(n289), .B(n290), .C(n291), .Z(n288) );
  GTECH_NOT U264 ( .A(n290), .Z(n286) );
  GTECH_NOT U265 ( .A(n292), .Z(n245) );
  GTECH_NAND2 U266 ( .A(I_a[5]), .B(I_b[3]), .Z(n292) );
  GTECH_NOT U267 ( .A(n241), .Z(n243) );
  GTECH_NAND2 U268 ( .A(I_a[6]), .B(I_b[2]), .Z(n241) );
  GTECH_XOR2 U269 ( .A(n293), .B(n250), .Z(n256) );
  GTECH_NOT U270 ( .A(n252), .Z(n250) );
  GTECH_OAI21 U271 ( .A(n285), .B(n294), .C(n295), .Z(n252) );
  GTECH_OAI21 U272 ( .A(n283), .B(n296), .C(n284), .Z(n295) );
  GTECH_NOT U273 ( .A(n296), .Z(n285) );
  GTECH_AND2 U274 ( .A(I_a[7]), .B(I_b[1]), .Z(n293) );
  GTECH_XOR2 U275 ( .A(n297), .B(n259), .Z(N147) );
  GTECH_ADD_ABC U276 ( .A(n298), .B(n299), .C(n300), .COUT(n259) );
  GTECH_XOR3 U277 ( .A(n301), .B(n302), .C(n303), .Z(n299) );
  GTECH_NOT U278 ( .A(n304), .Z(n302) );
  GTECH_OA21 U279 ( .A(n305), .B(n306), .C(n307), .Z(n298) );
  GTECH_XNOR4 U280 ( .A(n264), .B(n282), .C(n262), .D(n263), .Z(n297) );
  GTECH_ADD_ABC U281 ( .A(n301), .B(n308), .C(n303), .COUT(n263) );
  GTECH_NOT U282 ( .A(n309), .Z(n303) );
  GTECH_XOR3 U283 ( .A(n310), .B(n311), .C(n312), .Z(n308) );
  GTECH_XOR3 U284 ( .A(n270), .B(n229), .C(n228), .Z(n262) );
  GTECH_XOR2 U285 ( .A(n313), .B(n273), .Z(n228) );
  GTECH_NOT U286 ( .A(n314), .Z(n273) );
  GTECH_NAND2 U287 ( .A(I_b[7]), .B(I_a[0]), .Z(n314) );
  GTECH_NAND2 U288 ( .A(I_b[6]), .B(I_a[1]), .Z(n313) );
  GTECH_NOT U289 ( .A(n268), .Z(n229) );
  GTECH_XOR3 U290 ( .A(n277), .B(n279), .C(n278), .Z(n268) );
  GTECH_OAI21 U291 ( .A(n315), .B(n316), .C(n317), .Z(n278) );
  GTECH_NOT U292 ( .A(n318), .Z(n279) );
  GTECH_NAND2 U293 ( .A(I_b[5]), .B(I_a[2]), .Z(n318) );
  GTECH_NOT U294 ( .A(n275), .Z(n277) );
  GTECH_NAND2 U295 ( .A(I_b[4]), .B(I_a[3]), .Z(n275) );
  GTECH_NOT U296 ( .A(n319), .Z(n270) );
  GTECH_NAND3 U297 ( .A(I_a[0]), .B(n320), .C(I_b[6]), .Z(n319) );
  GTECH_NOT U298 ( .A(n321), .Z(n320) );
  GTECH_XOR3 U299 ( .A(n289), .B(n291), .C(n290), .Z(n282) );
  GTECH_OAI21 U300 ( .A(n322), .B(n323), .C(n324), .Z(n290) );
  GTECH_OAI21 U301 ( .A(n325), .B(n326), .C(n327), .Z(n324) );
  GTECH_NOT U302 ( .A(n326), .Z(n322) );
  GTECH_NOT U303 ( .A(n328), .Z(n291) );
  GTECH_NAND2 U304 ( .A(I_b[3]), .B(I_a[4]), .Z(n328) );
  GTECH_NOT U305 ( .A(n287), .Z(n289) );
  GTECH_NAND2 U306 ( .A(I_a[5]), .B(I_b[2]), .Z(n287) );
  GTECH_NOT U307 ( .A(n329), .Z(n264) );
  GTECH_XOR3 U308 ( .A(n283), .B(n284), .C(n296), .Z(n329) );
  GTECH_OAI21 U309 ( .A(n312), .B(n330), .C(n331), .Z(n296) );
  GTECH_OAI21 U310 ( .A(n310), .B(n332), .C(n311), .Z(n331) );
  GTECH_NOT U311 ( .A(n332), .Z(n312) );
  GTECH_NOT U312 ( .A(n333), .Z(n284) );
  GTECH_NAND2 U313 ( .A(I_a[6]), .B(I_b[1]), .Z(n333) );
  GTECH_NOT U314 ( .A(n294), .Z(n283) );
  GTECH_NAND2 U315 ( .A(I_a[7]), .B(I_b[0]), .Z(n294) );
  GTECH_XOR2 U316 ( .A(n334), .B(n335), .Z(N146) );
  GTECH_XNOR4 U317 ( .A(n309), .B(n301), .C(n304), .D(n300), .Z(n335) );
  GTECH_XOR2 U318 ( .A(n321), .B(n336), .Z(n300) );
  GTECH_AND2 U319 ( .A(I_b[6]), .B(I_a[0]), .Z(n336) );
  GTECH_XOR3 U320 ( .A(n337), .B(n338), .C(n317), .Z(n321) );
  GTECH_NAND3 U321 ( .A(I_b[4]), .B(I_a[1]), .C(n339), .Z(n317) );
  GTECH_NOT U322 ( .A(n316), .Z(n338) );
  GTECH_NAND2 U323 ( .A(I_b[5]), .B(I_a[1]), .Z(n316) );
  GTECH_NOT U324 ( .A(n315), .Z(n337) );
  GTECH_NAND2 U325 ( .A(I_b[4]), .B(I_a[2]), .Z(n315) );
  GTECH_XOR3 U326 ( .A(n310), .B(n311), .C(n332), .Z(n304) );
  GTECH_OAI21 U327 ( .A(n340), .B(n341), .C(n342), .Z(n332) );
  GTECH_OAI21 U328 ( .A(n343), .B(n344), .C(n345), .Z(n342) );
  GTECH_NOT U329 ( .A(n346), .Z(n311) );
  GTECH_NAND2 U330 ( .A(I_a[5]), .B(I_b[1]), .Z(n346) );
  GTECH_NOT U331 ( .A(n330), .Z(n310) );
  GTECH_NAND2 U332 ( .A(I_a[6]), .B(I_b[0]), .Z(n330) );
  GTECH_ADD_ABC U333 ( .A(n347), .B(n348), .C(n349), .COUT(n301) );
  GTECH_NOT U334 ( .A(n350), .Z(n349) );
  GTECH_XOR3 U335 ( .A(n343), .B(n345), .C(n340), .Z(n348) );
  GTECH_NOT U336 ( .A(n344), .Z(n340) );
  GTECH_XOR3 U337 ( .A(n325), .B(n327), .C(n326), .Z(n309) );
  GTECH_OAI21 U338 ( .A(n351), .B(n352), .C(n353), .Z(n326) );
  GTECH_OAI21 U339 ( .A(n354), .B(n355), .C(n356), .Z(n353) );
  GTECH_NOT U340 ( .A(n355), .Z(n351) );
  GTECH_NOT U341 ( .A(n357), .Z(n327) );
  GTECH_NAND2 U342 ( .A(I_b[3]), .B(I_a[3]), .Z(n357) );
  GTECH_NOT U343 ( .A(n323), .Z(n325) );
  GTECH_NAND2 U344 ( .A(I_b[2]), .B(I_a[4]), .Z(n323) );
  GTECH_OA21 U345 ( .A(n305), .B(n306), .C(n307), .Z(n334) );
  GTECH_OAI21 U346 ( .A(n358), .B(n359), .C(n360), .Z(n307) );
  GTECH_NOT U347 ( .A(n305), .Z(n359) );
  GTECH_XOR3 U348 ( .A(n360), .B(n306), .C(n305), .Z(N145) );
  GTECH_XOR2 U349 ( .A(n361), .B(n339), .Z(n305) );
  GTECH_NOT U350 ( .A(n362), .Z(n339) );
  GTECH_NAND2 U351 ( .A(I_b[5]), .B(I_a[0]), .Z(n362) );
  GTECH_NAND2 U352 ( .A(I_b[4]), .B(I_a[1]), .Z(n361) );
  GTECH_NOT U353 ( .A(n358), .Z(n306) );
  GTECH_XOR2 U354 ( .A(n363), .B(n347), .Z(n358) );
  GTECH_ADD_ABC U355 ( .A(n364), .B(n365), .C(n366), .COUT(n347) );
  GTECH_XOR3 U356 ( .A(n367), .B(n368), .C(n369), .Z(n365) );
  GTECH_OA21 U357 ( .A(n370), .B(n371), .C(n372), .Z(n364) );
  GTECH_XNOR4 U358 ( .A(n345), .B(n344), .C(n350), .D(n343), .Z(n363) );
  GTECH_NOT U359 ( .A(n341), .Z(n343) );
  GTECH_NAND2 U360 ( .A(I_a[5]), .B(I_b[0]), .Z(n341) );
  GTECH_XOR3 U361 ( .A(n354), .B(n356), .C(n355), .Z(n350) );
  GTECH_OAI21 U362 ( .A(n373), .B(n374), .C(n375), .Z(n355) );
  GTECH_NOT U363 ( .A(n376), .Z(n356) );
  GTECH_NAND2 U364 ( .A(I_b[3]), .B(I_a[2]), .Z(n376) );
  GTECH_NOT U365 ( .A(n352), .Z(n354) );
  GTECH_NAND2 U366 ( .A(I_b[2]), .B(I_a[3]), .Z(n352) );
  GTECH_OAI21 U367 ( .A(n369), .B(n377), .C(n378), .Z(n344) );
  GTECH_OAI21 U368 ( .A(n367), .B(n379), .C(n368), .Z(n378) );
  GTECH_NOT U369 ( .A(n377), .Z(n367) );
  GTECH_NOT U370 ( .A(n379), .Z(n369) );
  GTECH_NOT U371 ( .A(n380), .Z(n345) );
  GTECH_NAND2 U372 ( .A(I_a[4]), .B(I_b[1]), .Z(n380) );
  GTECH_NOT U373 ( .A(n381), .Z(n360) );
  GTECH_NAND3 U374 ( .A(I_a[0]), .B(n382), .C(I_b[4]), .Z(n381) );
  GTECH_XOR2 U375 ( .A(n383), .B(n382), .Z(N144) );
  GTECH_XOR2 U376 ( .A(n384), .B(n385), .Z(n382) );
  GTECH_XNOR4 U377 ( .A(n368), .B(n379), .C(n377), .D(n366), .Z(n385) );
  GTECH_XOR3 U378 ( .A(n386), .B(n387), .C(n375), .Z(n366) );
  GTECH_NAND3 U379 ( .A(I_b[2]), .B(I_a[1]), .C(n388), .Z(n375) );
  GTECH_NOT U380 ( .A(n374), .Z(n387) );
  GTECH_NAND2 U381 ( .A(I_b[3]), .B(I_a[1]), .Z(n374) );
  GTECH_NOT U382 ( .A(n373), .Z(n386) );
  GTECH_NAND2 U383 ( .A(I_b[2]), .B(I_a[2]), .Z(n373) );
  GTECH_NAND2 U384 ( .A(I_a[4]), .B(I_b[0]), .Z(n377) );
  GTECH_OAI21 U385 ( .A(n389), .B(n390), .C(n391), .Z(n379) );
  GTECH_OAI21 U386 ( .A(n392), .B(n393), .C(n394), .Z(n391) );
  GTECH_NOT U387 ( .A(n393), .Z(n389) );
  GTECH_NOT U388 ( .A(n395), .Z(n368) );
  GTECH_NAND2 U389 ( .A(I_a[3]), .B(I_b[1]), .Z(n395) );
  GTECH_OA21 U390 ( .A(n370), .B(n371), .C(n372), .Z(n384) );
  GTECH_OAI21 U391 ( .A(n396), .B(n397), .C(n398), .Z(n372) );
  GTECH_NOT U392 ( .A(n370), .Z(n397) );
  GTECH_AND2 U393 ( .A(I_b[4]), .B(I_a[0]), .Z(n383) );
  GTECH_XOR3 U394 ( .A(n398), .B(n371), .C(n370), .Z(N143) );
  GTECH_XOR2 U395 ( .A(n399), .B(n388), .Z(n370) );
  GTECH_NOT U396 ( .A(n400), .Z(n388) );
  GTECH_NAND2 U397 ( .A(I_b[3]), .B(I_a[0]), .Z(n400) );
  GTECH_NAND2 U398 ( .A(I_b[2]), .B(I_a[1]), .Z(n399) );
  GTECH_NOT U399 ( .A(n396), .Z(n371) );
  GTECH_XOR3 U400 ( .A(n392), .B(n394), .C(n393), .Z(n396) );
  GTECH_OAI21 U401 ( .A(n401), .B(n402), .C(n403), .Z(n393) );
  GTECH_NOT U402 ( .A(n404), .Z(n394) );
  GTECH_NAND2 U403 ( .A(I_b[1]), .B(I_a[2]), .Z(n404) );
  GTECH_NOT U404 ( .A(n390), .Z(n392) );
  GTECH_NAND2 U405 ( .A(I_b[0]), .B(I_a[3]), .Z(n390) );
  GTECH_NOT U406 ( .A(n405), .Z(n398) );
  GTECH_NAND3 U407 ( .A(I_a[0]), .B(n406), .C(I_b[2]), .Z(n405) );
  GTECH_XOR2 U408 ( .A(n407), .B(n406), .Z(N142) );
  GTECH_NOT U409 ( .A(n408), .Z(n406) );
  GTECH_XOR3 U410 ( .A(n409), .B(n410), .C(n403), .Z(n408) );
  GTECH_NAND3 U411 ( .A(n411), .B(I_b[0]), .C(I_a[1]), .Z(n403) );
  GTECH_NOT U412 ( .A(n401), .Z(n410) );
  GTECH_NAND2 U413 ( .A(I_a[1]), .B(I_b[1]), .Z(n401) );
  GTECH_NOT U414 ( .A(n402), .Z(n409) );
  GTECH_NAND2 U415 ( .A(I_b[0]), .B(I_a[2]), .Z(n402) );
  GTECH_AND2 U416 ( .A(I_b[2]), .B(I_a[0]), .Z(n407) );
  GTECH_XOR2 U417 ( .A(n411), .B(n412), .Z(N141) );
  GTECH_AND2 U418 ( .A(I_a[1]), .B(I_b[0]), .Z(n412) );
  GTECH_NOT U419 ( .A(n413), .Z(n411) );
  GTECH_NAND2 U420 ( .A(I_a[0]), .B(I_b[1]), .Z(n413) );
  GTECH_AND2 U421 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

