
module fraction_multiplier4 ( CLK, St, Mplier, Mcand, Product, Done );
  input [3:0] Mplier;
  input [3:0] Mcand;
  output [6:0] Product;
  input CLK, St;
  output Done;
  wire   N40, N41, N42, N44, N46, N48, N50, N52, N54, N56, N57, N58, N63, n12,
         n14, n15, n16, n17, n18, n19, n73, n81, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139;
  wire   [2:0] State;

  GTECH_FD2 State_reg_0_ ( .D(N40), .CP(CLK), .CD(n81), .Q(State[0]), .QN(n85)
         );
  GTECH_FD2 State_reg_2_ ( .D(N42), .CP(CLK), .CD(n81), .Q(State[2]), .QN(n87)
         );
  GTECH_FD2 State_reg_1_ ( .D(N41), .CP(CLK), .CD(n81), .Q(State[1]), .QN(n86)
         );
  GTECH_FJK1S B_reg_0_ ( .J(n73), .K(n73), .TI(N52), .TE(N57), .CP(CLK), .Q(
        Product[0]), .QN(n12) );
  GTECH_FJK1S A_reg_3_ ( .J(n73), .K(n73), .TI(N50), .TE(N63), .CP(CLK), .QN(
        n84) );
  GTECH_FJK1S A_reg_0_ ( .J(n73), .K(n73), .TI(N44), .TE(N57), .CP(CLK), .Q(
        Product[4]), .QN(n14) );
  GTECH_FJK1S A_reg_1_ ( .J(n73), .K(n73), .TI(N46), .TE(N57), .CP(CLK), .Q(
        Product[5]), .QN(n15) );
  GTECH_FJK1S A_reg_2_ ( .J(n73), .K(n73), .TI(N48), .TE(N57), .CP(CLK), .Q(
        Product[6]), .QN(n16) );
  GTECH_FJK1S B_reg_3_ ( .J(n73), .K(n73), .TI(N58), .TE(N57), .CP(CLK), .Q(
        Product[3]), .QN(n17) );
  GTECH_FJK1S B_reg_2_ ( .J(n73), .K(n73), .TI(N56), .TE(N57), .CP(CLK), .Q(
        Product[2]), .QN(n18) );
  GTECH_FJK1S B_reg_1_ ( .J(n73), .K(n73), .TI(N54), .TE(N57), .CP(CLK), .Q(
        Product[1]), .QN(n19) );
  GTECH_ONE U81 ( .Z(n81) );
  GTECH_ZERO U82 ( .Z(n73) );
  GTECH_AND2 U83 ( .A(n88), .B(N57), .Z(N63) );
  GTECH_NOT U84 ( .A(n89), .Z(N58) );
  GTECH_AOI222 U85 ( .A(Mplier[3]), .B(n90), .C(n91), .D(n92), .E(n93), .F(n94), .Z(n89) );
  GTECH_OAI21 U86 ( .A(Mcand[0]), .B(n95), .C(n88), .Z(n93) );
  GTECH_NOR2 U87 ( .A(n95), .B(n12), .Z(n91) );
  GTECH_OAI21 U88 ( .A(n96), .B(n97), .C(n95), .Z(N57) );
  GTECH_OAI2N2 U89 ( .A(n17), .B(n95), .C(Mplier[2]), .D(n90), .Z(N56) );
  GTECH_OAI2N2 U90 ( .A(n18), .B(n95), .C(Mplier[1]), .D(n90), .Z(N54) );
  GTECH_OAI2N2 U91 ( .A(n19), .B(n95), .C(Mplier[0]), .D(n90), .Z(N52) );
  GTECH_MUX2 U92 ( .A(n98), .B(n99), .S(Mcand[3]), .Z(N50) );
  GTECH_MUX2 U93 ( .A(n100), .B(n101), .S(n84), .Z(N48) );
  GTECH_MUX2 U94 ( .A(n102), .B(n103), .S(Mcand[3]), .Z(n101) );
  GTECH_OR_NOT U95 ( .A(n104), .B(n88), .Z(n100) );
  GTECH_MUX2 U96 ( .A(n103), .B(n102), .S(Mcand[3]), .Z(n104) );
  GTECH_OAI2N2 U97 ( .A(n105), .B(n106), .C(n107), .D(n108), .Z(n102) );
  GTECH_OAI2N2 U98 ( .A(n107), .B(n109), .C(n110), .D(n105), .Z(n103) );
  GTECH_OA21 U99 ( .A(n111), .B(n112), .C(n113), .Z(n105) );
  GTECH_AO21 U100 ( .A(n112), .B(n111), .C(n16), .Z(n113) );
  GTECH_NOT U101 ( .A(Mcand[2]), .Z(n112) );
  GTECH_ADD_ABC U102 ( .A(Mcand[2]), .B(n114), .C(n16), .COUT(n107) );
  GTECH_MUX2 U103 ( .A(n115), .B(n116), .S(n16), .Z(N46) );
  GTECH_NOT U104 ( .A(n117), .Z(n116) );
  GTECH_MUX2 U105 ( .A(n118), .B(n119), .S(Mcand[2]), .Z(n117) );
  GTECH_NAND2 U106 ( .A(n120), .B(n88), .Z(n115) );
  GTECH_MUX2 U107 ( .A(n119), .B(n118), .S(Mcand[2]), .Z(n120) );
  GTECH_AOI2N2 U108 ( .A(n114), .B(n108), .C(n111), .D(n106), .Z(n118) );
  GTECH_AOI2N2 U109 ( .A(n111), .B(n110), .C(n114), .D(n109), .Z(n119) );
  GTECH_ADD_ABC U110 ( .A(Mcand[1]), .B(n92), .C(n15), .COUT(n114) );
  GTECH_OA21 U111 ( .A(n15), .B(n121), .C(n122), .Z(n111) );
  GTECH_OR3 U112 ( .A(n123), .B(n14), .C(n124), .Z(n122) );
  GTECH_NAND2 U113 ( .A(n125), .B(n126), .Z(N44) );
  GTECH_MUX2 U114 ( .A(n127), .B(n128), .S(n15), .Z(n126) );
  GTECH_OR_NOT U115 ( .A(n121), .B(n129), .Z(n128) );
  GTECH_AND_NOT U116 ( .A(n88), .B(n130), .Z(n127) );
  GTECH_MUX2 U117 ( .A(n131), .B(n129), .S(n121), .Z(n130) );
  GTECH_OAI21 U118 ( .A(n92), .B(n109), .C(n132), .Z(n129) );
  GTECH_AO21 U119 ( .A(n94), .B(Mcand[0]), .C(n106), .Z(n132) );
  GTECH_NOT U120 ( .A(n108), .Z(n109) );
  GTECH_AND_NOT U121 ( .A(Mcand[0]), .B(n94), .Z(n92) );
  GTECH_NOT U122 ( .A(n14), .Z(n94) );
  GTECH_AND_NOT U123 ( .A(n133), .B(n124), .Z(n131) );
  GTECH_NOT U124 ( .A(Mcand[0]), .Z(n124) );
  GTECH_OR_NOT U125 ( .A(n95), .B(n12), .Z(n88) );
  GTECH_NOR2 U126 ( .A(n98), .B(n99), .Z(n95) );
  GTECH_NAND3 U127 ( .A(Mcand[0]), .B(n133), .C(n123), .Z(n125) );
  GTECH_AND2 U128 ( .A(n15), .B(n121), .Z(n123) );
  GTECH_NOT U129 ( .A(Mcand[1]), .Z(n121) );
  GTECH_MUX2 U130 ( .A(n110), .B(n108), .S(n14), .Z(n133) );
  GTECH_NOR2 U131 ( .A(n134), .B(n12), .Z(n108) );
  GTECH_NOT U132 ( .A(n98), .Z(n134) );
  GTECH_NOT U133 ( .A(n106), .Z(n110) );
  GTECH_OR_NOT U134 ( .A(n12), .B(n99), .Z(n106) );
  GTECH_OR_NOT U135 ( .A(n98), .B(n135), .Z(N42) );
  GTECH_NAND3 U136 ( .A(n136), .B(n137), .C(n99), .Z(n135) );
  GTECH_OA21 U137 ( .A(n85), .B(n86), .C(n99), .Z(N41) );
  GTECH_OAI21 U138 ( .A(n96), .B(n97), .C(n138), .Z(N40) );
  GTECH_AOI21 U139 ( .A(n85), .B(n99), .C(n98), .Z(n138) );
  GTECH_NOR3 U140 ( .A(n136), .B(n87), .C(n137), .Z(n98) );
  GTECH_AOI21 U141 ( .A(n85), .B(n86), .C(n139), .Z(n99) );
  GTECH_NOT U142 ( .A(St), .Z(n97) );
  GTECH_NOT U143 ( .A(n90), .Z(n96) );
  GTECH_NOR3 U144 ( .A(n137), .B(n136), .C(n139), .Z(n90) );
  GTECH_NOT U145 ( .A(n87), .Z(n139) );
  GTECH_NOT U146 ( .A(n85), .Z(n136) );
  GTECH_NOR3 U147 ( .A(n85), .B(n87), .C(n137), .Z(Done) );
  GTECH_NOT U148 ( .A(n86), .Z(n137) );
endmodule

