
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_OAI21 U75 ( .A(n83), .B(n84), .C(n85), .Z(N155) );
  GTECH_OA22 U76 ( .A(n86), .B(n87), .C(n88), .D(n89), .Z(n85) );
  GTECH_NOT U77 ( .A(n90), .Z(n87) );
  GTECH_XOR2 U78 ( .A(n91), .B(n92), .Z(N154) );
  GTECH_NOT U79 ( .A(n83), .Z(n92) );
  GTECH_XOR2 U80 ( .A(n90), .B(n86), .Z(n83) );
  GTECH_AOI2N2 U81 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n86) );
  GTECH_NAND2 U82 ( .A(n95), .B(n96), .Z(n94) );
  GTECH_XOR2 U83 ( .A(n89), .B(n88), .Z(n90) );
  GTECH_AND2 U84 ( .A(n97), .B(n98), .Z(n88) );
  GTECH_OR_NOT U85 ( .A(n99), .B(n100), .Z(n98) );
  GTECH_OAI21 U86 ( .A(n101), .B(n100), .C(n102), .Z(n97) );
  GTECH_NAND2 U87 ( .A(I_b[7]), .B(I_a[7]), .Z(n89) );
  GTECH_NOT U88 ( .A(n84), .Z(n91) );
  GTECH_NAND2 U89 ( .A(n103), .B(n104), .Z(n84) );
  GTECH_XOR2 U90 ( .A(n104), .B(n103), .Z(N153) );
  GTECH_NOT U91 ( .A(n105), .Z(n103) );
  GTECH_XOR3 U92 ( .A(n106), .B(n95), .C(n93), .Z(n105) );
  GTECH_XOR3 U93 ( .A(n101), .B(n102), .C(n100), .Z(n93) );
  GTECH_OAI21 U94 ( .A(n107), .B(n108), .C(n109), .Z(n100) );
  GTECH_OAI21 U95 ( .A(n110), .B(n111), .C(n112), .Z(n109) );
  GTECH_NOT U96 ( .A(n111), .Z(n107) );
  GTECH_NOT U97 ( .A(n113), .Z(n102) );
  GTECH_NAND2 U98 ( .A(I_b[7]), .B(I_a[6]), .Z(n113) );
  GTECH_NOT U99 ( .A(n99), .Z(n101) );
  GTECH_NAND2 U100 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U101 ( .A(n114), .B(n115), .C(n116), .COUT(n95) );
  GTECH_NOT U102 ( .A(n117), .Z(n116) );
  GTECH_XOR2 U103 ( .A(n118), .B(n119), .Z(n115) );
  GTECH_AND2 U104 ( .A(I_a[7]), .B(I_b[5]), .Z(n119) );
  GTECH_NOT U105 ( .A(n96), .Z(n106) );
  GTECH_NAND2 U106 ( .A(I_a[7]), .B(n120), .Z(n96) );
  GTECH_NOT U107 ( .A(n121), .Z(n104) );
  GTECH_NAND2 U108 ( .A(n122), .B(n123), .Z(n121) );
  GTECH_NOT U109 ( .A(n124), .Z(n123) );
  GTECH_XOR2 U110 ( .A(n124), .B(n125), .Z(N152) );
  GTECH_NOT U111 ( .A(n122), .Z(n125) );
  GTECH_XOR4 U112 ( .A(n126), .B(n118), .C(n114), .D(n117), .Z(n122) );
  GTECH_XOR3 U113 ( .A(n110), .B(n112), .C(n111), .Z(n117) );
  GTECH_OAI21 U114 ( .A(n127), .B(n128), .C(n129), .Z(n111) );
  GTECH_OAI21 U115 ( .A(n130), .B(n131), .C(n132), .Z(n129) );
  GTECH_NOT U116 ( .A(n131), .Z(n127) );
  GTECH_NOT U117 ( .A(n133), .Z(n112) );
  GTECH_NAND2 U118 ( .A(I_b[7]), .B(I_a[5]), .Z(n133) );
  GTECH_NOT U119 ( .A(n108), .Z(n110) );
  GTECH_NAND2 U120 ( .A(I_b[6]), .B(I_a[6]), .Z(n108) );
  GTECH_ADD_ABC U121 ( .A(n134), .B(n135), .C(n136), .COUT(n114) );
  GTECH_NOT U122 ( .A(n137), .Z(n136) );
  GTECH_XOR3 U123 ( .A(n138), .B(n139), .C(n140), .Z(n135) );
  GTECH_NOT U124 ( .A(n120), .Z(n118) );
  GTECH_OAI21 U125 ( .A(n140), .B(n141), .C(n142), .Z(n120) );
  GTECH_OAI21 U126 ( .A(n138), .B(n143), .C(n139), .Z(n142) );
  GTECH_NOT U127 ( .A(n141), .Z(n138) );
  GTECH_NOT U128 ( .A(n143), .Z(n140) );
  GTECH_AND2 U129 ( .A(I_a[7]), .B(I_b[5]), .Z(n126) );
  GTECH_ADD_ABC U130 ( .A(n144), .B(n145), .C(n146), .COUT(n124) );
  GTECH_NOT U131 ( .A(n147), .Z(n146) );
  GTECH_OA22 U132 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n145) );
  GTECH_OA21 U133 ( .A(n152), .B(n153), .C(n154), .Z(n144) );
  GTECH_XOR3 U134 ( .A(n155), .B(n147), .C(n156), .Z(N151) );
  GTECH_OA21 U135 ( .A(n152), .B(n153), .C(n154), .Z(n156) );
  GTECH_OAI21 U136 ( .A(n157), .B(n158), .C(n159), .Z(n154) );
  GTECH_XOR2 U137 ( .A(n160), .B(n134), .Z(n147) );
  GTECH_ADD_ABC U138 ( .A(n161), .B(n162), .C(n163), .COUT(n134) );
  GTECH_NOT U139 ( .A(n164), .Z(n163) );
  GTECH_XOR3 U140 ( .A(n165), .B(n166), .C(n167), .Z(n162) );
  GTECH_XOR4 U141 ( .A(n139), .B(n143), .C(n141), .D(n137), .Z(n160) );
  GTECH_XOR3 U142 ( .A(n130), .B(n132), .C(n131), .Z(n137) );
  GTECH_OAI21 U143 ( .A(n168), .B(n169), .C(n170), .Z(n131) );
  GTECH_OAI21 U144 ( .A(n171), .B(n172), .C(n173), .Z(n170) );
  GTECH_NOT U145 ( .A(n172), .Z(n168) );
  GTECH_NOT U146 ( .A(n174), .Z(n132) );
  GTECH_NAND2 U147 ( .A(I_b[7]), .B(I_a[4]), .Z(n174) );
  GTECH_NOT U148 ( .A(n128), .Z(n130) );
  GTECH_NAND2 U149 ( .A(I_b[6]), .B(I_a[5]), .Z(n128) );
  GTECH_NAND2 U150 ( .A(I_a[7]), .B(I_b[4]), .Z(n141) );
  GTECH_OAI21 U151 ( .A(n167), .B(n175), .C(n176), .Z(n143) );
  GTECH_OAI21 U152 ( .A(n165), .B(n177), .C(n166), .Z(n176) );
  GTECH_NOT U153 ( .A(n175), .Z(n165) );
  GTECH_NOT U154 ( .A(n177), .Z(n167) );
  GTECH_NOT U155 ( .A(n178), .Z(n139) );
  GTECH_NAND2 U156 ( .A(I_a[6]), .B(I_b[5]), .Z(n178) );
  GTECH_OA22 U157 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n155) );
  GTECH_NOT U158 ( .A(n179), .Z(n151) );
  GTECH_NOT U159 ( .A(I_a[7]), .Z(n149) );
  GTECH_XOR3 U160 ( .A(n152), .B(n157), .C(n180), .Z(N150) );
  GTECH_NOT U161 ( .A(n159), .Z(n180) );
  GTECH_XOR2 U162 ( .A(n181), .B(n161), .Z(n159) );
  GTECH_ADD_ABC U163 ( .A(n182), .B(n183), .C(n184), .COUT(n161) );
  GTECH_NOT U164 ( .A(n185), .Z(n184) );
  GTECH_XOR3 U165 ( .A(n186), .B(n187), .C(n188), .Z(n183) );
  GTECH_XOR4 U166 ( .A(n166), .B(n177), .C(n175), .D(n164), .Z(n181) );
  GTECH_XOR3 U167 ( .A(n171), .B(n173), .C(n172), .Z(n164) );
  GTECH_OAI21 U168 ( .A(n189), .B(n190), .C(n191), .Z(n172) );
  GTECH_OAI21 U169 ( .A(n192), .B(n193), .C(n194), .Z(n191) );
  GTECH_NOT U170 ( .A(n193), .Z(n189) );
  GTECH_NOT U171 ( .A(n195), .Z(n173) );
  GTECH_NAND2 U172 ( .A(I_b[7]), .B(I_a[3]), .Z(n195) );
  GTECH_NOT U173 ( .A(n169), .Z(n171) );
  GTECH_NAND2 U174 ( .A(I_b[6]), .B(I_a[4]), .Z(n169) );
  GTECH_NAND2 U175 ( .A(I_a[6]), .B(I_b[4]), .Z(n175) );
  GTECH_OAI21 U176 ( .A(n188), .B(n196), .C(n197), .Z(n177) );
  GTECH_OAI21 U177 ( .A(n186), .B(n198), .C(n187), .Z(n197) );
  GTECH_NOT U178 ( .A(n196), .Z(n186) );
  GTECH_NOT U179 ( .A(n198), .Z(n188) );
  GTECH_NOT U180 ( .A(n199), .Z(n166) );
  GTECH_NAND2 U181 ( .A(I_a[5]), .B(I_b[5]), .Z(n199) );
  GTECH_NOT U182 ( .A(n153), .Z(n157) );
  GTECH_XOR2 U183 ( .A(n179), .B(n150), .Z(n153) );
  GTECH_AOI2N2 U184 ( .A(n200), .B(n201), .C(n202), .D(n203), .Z(n150) );
  GTECH_NAND2 U185 ( .A(n202), .B(n203), .Z(n201) );
  GTECH_XOR2 U186 ( .A(n204), .B(n148), .Z(n179) );
  GTECH_AND2 U187 ( .A(n205), .B(n206), .Z(n148) );
  GTECH_OR_NOT U188 ( .A(n207), .B(n208), .Z(n206) );
  GTECH_OAI21 U189 ( .A(n209), .B(n208), .C(n210), .Z(n205) );
  GTECH_NAND2 U190 ( .A(I_a[7]), .B(I_b[3]), .Z(n204) );
  GTECH_NOT U191 ( .A(n158), .Z(n152) );
  GTECH_OAI21 U192 ( .A(n211), .B(n212), .C(n213), .Z(n158) );
  GTECH_OAI21 U193 ( .A(n214), .B(n215), .C(n216), .Z(n213) );
  GTECH_NOT U194 ( .A(n211), .Z(n215) );
  GTECH_XOR3 U195 ( .A(n211), .B(n214), .C(n217), .Z(N149) );
  GTECH_NOT U196 ( .A(n216), .Z(n217) );
  GTECH_XOR2 U197 ( .A(n218), .B(n182), .Z(n216) );
  GTECH_ADD_ABC U198 ( .A(n219), .B(n220), .C(n221), .COUT(n182) );
  GTECH_XOR3 U199 ( .A(n222), .B(n223), .C(n224), .Z(n220) );
  GTECH_OA21 U200 ( .A(n225), .B(n226), .C(n227), .Z(n219) );
  GTECH_XOR4 U201 ( .A(n187), .B(n198), .C(n196), .D(n185), .Z(n218) );
  GTECH_XOR3 U202 ( .A(n192), .B(n194), .C(n193), .Z(n185) );
  GTECH_OAI21 U203 ( .A(n228), .B(n229), .C(n230), .Z(n193) );
  GTECH_NOT U204 ( .A(n231), .Z(n194) );
  GTECH_NAND2 U205 ( .A(I_b[7]), .B(I_a[2]), .Z(n231) );
  GTECH_NOT U206 ( .A(n190), .Z(n192) );
  GTECH_NAND2 U207 ( .A(I_b[6]), .B(I_a[3]), .Z(n190) );
  GTECH_NAND2 U208 ( .A(I_a[5]), .B(I_b[4]), .Z(n196) );
  GTECH_OAI21 U209 ( .A(n224), .B(n232), .C(n233), .Z(n198) );
  GTECH_OAI21 U210 ( .A(n222), .B(n234), .C(n223), .Z(n233) );
  GTECH_NOT U211 ( .A(n232), .Z(n222) );
  GTECH_NOT U212 ( .A(n234), .Z(n224) );
  GTECH_NOT U213 ( .A(n235), .Z(n187) );
  GTECH_NAND2 U214 ( .A(I_b[5]), .B(I_a[4]), .Z(n235) );
  GTECH_NOT U215 ( .A(n212), .Z(n214) );
  GTECH_XOR3 U216 ( .A(n236), .B(n202), .C(n200), .Z(n212) );
  GTECH_XOR3 U217 ( .A(n209), .B(n210), .C(n208), .Z(n200) );
  GTECH_OAI21 U218 ( .A(n237), .B(n238), .C(n239), .Z(n208) );
  GTECH_OAI21 U219 ( .A(n240), .B(n241), .C(n242), .Z(n239) );
  GTECH_NOT U220 ( .A(n241), .Z(n237) );
  GTECH_NOT U221 ( .A(n243), .Z(n210) );
  GTECH_NAND2 U222 ( .A(I_a[6]), .B(I_b[3]), .Z(n243) );
  GTECH_NOT U223 ( .A(n207), .Z(n209) );
  GTECH_NAND2 U224 ( .A(I_a[7]), .B(I_b[2]), .Z(n207) );
  GTECH_ADD_ABC U225 ( .A(n244), .B(n245), .C(n246), .COUT(n202) );
  GTECH_XOR2 U226 ( .A(n247), .B(n248), .Z(n245) );
  GTECH_AND2 U227 ( .A(I_a[7]), .B(I_b[1]), .Z(n248) );
  GTECH_NOT U228 ( .A(n203), .Z(n236) );
  GTECH_NAND2 U229 ( .A(I_a[7]), .B(n249), .Z(n203) );
  GTECH_ADD_ABC U230 ( .A(n250), .B(n251), .C(n252), .COUT(n211) );
  GTECH_XOR3 U231 ( .A(n244), .B(n253), .C(n246), .Z(n251) );
  GTECH_NOT U232 ( .A(n254), .Z(n246) );
  GTECH_XOR2 U233 ( .A(n250), .B(n255), .Z(N148) );
  GTECH_XOR4 U234 ( .A(n253), .B(n254), .C(n252), .D(n244), .Z(n255) );
  GTECH_ADD_ABC U235 ( .A(n256), .B(n257), .C(n258), .COUT(n244) );
  GTECH_XOR3 U236 ( .A(n259), .B(n260), .C(n261), .Z(n257) );
  GTECH_XOR2 U237 ( .A(n262), .B(n263), .Z(n252) );
  GTECH_OA21 U238 ( .A(n225), .B(n226), .C(n227), .Z(n263) );
  GTECH_OAI21 U239 ( .A(n264), .B(n265), .C(n266), .Z(n227) );
  GTECH_NOT U240 ( .A(n225), .Z(n265) );
  GTECH_XOR4 U241 ( .A(n223), .B(n234), .C(n232), .D(n221), .Z(n262) );
  GTECH_XOR3 U242 ( .A(n267), .B(n268), .C(n230), .Z(n221) );
  GTECH_NAND3 U243 ( .A(I_b[6]), .B(I_a[1]), .C(n269), .Z(n230) );
  GTECH_NOT U244 ( .A(n229), .Z(n268) );
  GTECH_NAND2 U245 ( .A(I_b[7]), .B(I_a[1]), .Z(n229) );
  GTECH_NOT U246 ( .A(n228), .Z(n267) );
  GTECH_NAND2 U247 ( .A(I_b[6]), .B(I_a[2]), .Z(n228) );
  GTECH_NAND2 U248 ( .A(I_b[4]), .B(I_a[4]), .Z(n232) );
  GTECH_OAI21 U249 ( .A(n270), .B(n271), .C(n272), .Z(n234) );
  GTECH_OAI21 U250 ( .A(n273), .B(n274), .C(n275), .Z(n272) );
  GTECH_NOT U251 ( .A(n274), .Z(n270) );
  GTECH_NOT U252 ( .A(n276), .Z(n223) );
  GTECH_NAND2 U253 ( .A(I_b[5]), .B(I_a[3]), .Z(n276) );
  GTECH_XOR3 U254 ( .A(n240), .B(n242), .C(n241), .Z(n254) );
  GTECH_OAI21 U255 ( .A(n277), .B(n278), .C(n279), .Z(n241) );
  GTECH_OAI21 U256 ( .A(n280), .B(n281), .C(n282), .Z(n279) );
  GTECH_NOT U257 ( .A(n281), .Z(n277) );
  GTECH_NOT U258 ( .A(n283), .Z(n242) );
  GTECH_NAND2 U259 ( .A(I_a[5]), .B(I_b[3]), .Z(n283) );
  GTECH_NOT U260 ( .A(n238), .Z(n240) );
  GTECH_NAND2 U261 ( .A(I_a[6]), .B(I_b[2]), .Z(n238) );
  GTECH_XOR2 U262 ( .A(n284), .B(n247), .Z(n253) );
  GTECH_NOT U263 ( .A(n249), .Z(n247) );
  GTECH_OAI21 U264 ( .A(n261), .B(n285), .C(n286), .Z(n249) );
  GTECH_OAI21 U265 ( .A(n259), .B(n287), .C(n260), .Z(n286) );
  GTECH_NOT U266 ( .A(n287), .Z(n261) );
  GTECH_AND2 U267 ( .A(I_a[7]), .B(I_b[1]), .Z(n284) );
  GTECH_ADD_ABC U268 ( .A(n288), .B(n289), .C(n290), .COUT(n250) );
  GTECH_NOT U269 ( .A(n291), .Z(n290) );
  GTECH_XOR3 U270 ( .A(n256), .B(n292), .C(n258), .Z(n289) );
  GTECH_NOT U271 ( .A(n293), .Z(n258) );
  GTECH_NOT U272 ( .A(n294), .Z(n292) );
  GTECH_XOR2 U273 ( .A(n295), .B(n288), .Z(N147) );
  GTECH_ADD_ABC U274 ( .A(n296), .B(n297), .C(n298), .COUT(n288) );
  GTECH_XOR3 U275 ( .A(n299), .B(n300), .C(n301), .Z(n297) );
  GTECH_OA21 U276 ( .A(n302), .B(n303), .C(n304), .Z(n296) );
  GTECH_XOR4 U277 ( .A(n293), .B(n256), .C(n294), .D(n291), .Z(n295) );
  GTECH_XOR3 U278 ( .A(n266), .B(n226), .C(n225), .Z(n291) );
  GTECH_XOR2 U279 ( .A(n305), .B(n269), .Z(n225) );
  GTECH_NOT U280 ( .A(n306), .Z(n269) );
  GTECH_NAND2 U281 ( .A(I_b[7]), .B(I_a[0]), .Z(n306) );
  GTECH_NAND2 U282 ( .A(I_b[6]), .B(I_a[1]), .Z(n305) );
  GTECH_NOT U283 ( .A(n264), .Z(n226) );
  GTECH_XOR3 U284 ( .A(n273), .B(n275), .C(n274), .Z(n264) );
  GTECH_OAI21 U285 ( .A(n307), .B(n308), .C(n309), .Z(n274) );
  GTECH_NOT U286 ( .A(n310), .Z(n275) );
  GTECH_NAND2 U287 ( .A(I_b[5]), .B(I_a[2]), .Z(n310) );
  GTECH_NOT U288 ( .A(n271), .Z(n273) );
  GTECH_NAND2 U289 ( .A(I_b[4]), .B(I_a[3]), .Z(n271) );
  GTECH_NOT U290 ( .A(n311), .Z(n266) );
  GTECH_NAND3 U291 ( .A(I_a[0]), .B(n312), .C(I_b[6]), .Z(n311) );
  GTECH_NOT U292 ( .A(n313), .Z(n312) );
  GTECH_XOR3 U293 ( .A(n259), .B(n260), .C(n287), .Z(n294) );
  GTECH_OAI21 U294 ( .A(n314), .B(n315), .C(n316), .Z(n287) );
  GTECH_OAI21 U295 ( .A(n317), .B(n318), .C(n319), .Z(n316) );
  GTECH_NOT U296 ( .A(n320), .Z(n260) );
  GTECH_NAND2 U297 ( .A(I_a[6]), .B(I_b[1]), .Z(n320) );
  GTECH_NOT U298 ( .A(n285), .Z(n259) );
  GTECH_NAND2 U299 ( .A(I_a[7]), .B(I_b[0]), .Z(n285) );
  GTECH_ADD_ABC U300 ( .A(n299), .B(n321), .C(n301), .COUT(n256) );
  GTECH_NOT U301 ( .A(n322), .Z(n301) );
  GTECH_XOR3 U302 ( .A(n317), .B(n319), .C(n314), .Z(n321) );
  GTECH_NOT U303 ( .A(n318), .Z(n314) );
  GTECH_XOR3 U304 ( .A(n280), .B(n282), .C(n281), .Z(n293) );
  GTECH_OAI21 U305 ( .A(n323), .B(n324), .C(n325), .Z(n281) );
  GTECH_OAI21 U306 ( .A(n326), .B(n327), .C(n328), .Z(n325) );
  GTECH_NOT U307 ( .A(n327), .Z(n323) );
  GTECH_NOT U308 ( .A(n329), .Z(n282) );
  GTECH_NAND2 U309 ( .A(I_b[3]), .B(I_a[4]), .Z(n329) );
  GTECH_NOT U310 ( .A(n278), .Z(n280) );
  GTECH_NAND2 U311 ( .A(I_a[5]), .B(I_b[2]), .Z(n278) );
  GTECH_XOR2 U312 ( .A(n330), .B(n331), .Z(N146) );
  GTECH_XOR4 U313 ( .A(n300), .B(n322), .C(n298), .D(n299), .Z(n331) );
  GTECH_ADD_ABC U314 ( .A(n332), .B(n333), .C(n334), .COUT(n299) );
  GTECH_NOT U315 ( .A(n335), .Z(n334) );
  GTECH_XOR3 U316 ( .A(n336), .B(n337), .C(n338), .Z(n333) );
  GTECH_XOR2 U317 ( .A(n313), .B(n339), .Z(n298) );
  GTECH_AND2 U318 ( .A(I_b[6]), .B(I_a[0]), .Z(n339) );
  GTECH_XOR3 U319 ( .A(n340), .B(n341), .C(n309), .Z(n313) );
  GTECH_NAND3 U320 ( .A(I_b[4]), .B(I_a[1]), .C(n342), .Z(n309) );
  GTECH_NOT U321 ( .A(n308), .Z(n341) );
  GTECH_NAND2 U322 ( .A(I_b[5]), .B(I_a[1]), .Z(n308) );
  GTECH_NOT U323 ( .A(n307), .Z(n340) );
  GTECH_NAND2 U324 ( .A(I_b[4]), .B(I_a[2]), .Z(n307) );
  GTECH_XOR3 U325 ( .A(n326), .B(n328), .C(n327), .Z(n322) );
  GTECH_OAI21 U326 ( .A(n343), .B(n344), .C(n345), .Z(n327) );
  GTECH_OAI21 U327 ( .A(n346), .B(n347), .C(n348), .Z(n345) );
  GTECH_NOT U328 ( .A(n347), .Z(n343) );
  GTECH_NOT U329 ( .A(n349), .Z(n328) );
  GTECH_NAND2 U330 ( .A(I_b[3]), .B(I_a[3]), .Z(n349) );
  GTECH_NOT U331 ( .A(n324), .Z(n326) );
  GTECH_NAND2 U332 ( .A(I_b[2]), .B(I_a[4]), .Z(n324) );
  GTECH_NOT U333 ( .A(n350), .Z(n300) );
  GTECH_XOR3 U334 ( .A(n317), .B(n319), .C(n318), .Z(n350) );
  GTECH_OAI21 U335 ( .A(n338), .B(n351), .C(n352), .Z(n318) );
  GTECH_OAI21 U336 ( .A(n336), .B(n353), .C(n337), .Z(n352) );
  GTECH_NOT U337 ( .A(n351), .Z(n336) );
  GTECH_NOT U338 ( .A(n353), .Z(n338) );
  GTECH_NOT U339 ( .A(n354), .Z(n319) );
  GTECH_NAND2 U340 ( .A(I_a[5]), .B(I_b[1]), .Z(n354) );
  GTECH_NOT U341 ( .A(n315), .Z(n317) );
  GTECH_NAND2 U342 ( .A(I_a[6]), .B(I_b[0]), .Z(n315) );
  GTECH_OA21 U343 ( .A(n302), .B(n303), .C(n304), .Z(n330) );
  GTECH_OAI21 U344 ( .A(n355), .B(n356), .C(n357), .Z(n304) );
  GTECH_NOT U345 ( .A(n302), .Z(n356) );
  GTECH_XOR3 U346 ( .A(n357), .B(n303), .C(n302), .Z(N145) );
  GTECH_XOR2 U347 ( .A(n358), .B(n342), .Z(n302) );
  GTECH_NOT U348 ( .A(n359), .Z(n342) );
  GTECH_NAND2 U349 ( .A(I_b[5]), .B(I_a[0]), .Z(n359) );
  GTECH_NAND2 U350 ( .A(I_b[4]), .B(I_a[1]), .Z(n358) );
  GTECH_NOT U351 ( .A(n355), .Z(n303) );
  GTECH_XOR2 U352 ( .A(n360), .B(n332), .Z(n355) );
  GTECH_ADD_ABC U353 ( .A(n361), .B(n362), .C(n363), .COUT(n332) );
  GTECH_XOR3 U354 ( .A(n364), .B(n365), .C(n366), .Z(n362) );
  GTECH_OA21 U355 ( .A(n367), .B(n368), .C(n369), .Z(n361) );
  GTECH_XOR4 U356 ( .A(n337), .B(n353), .C(n351), .D(n335), .Z(n360) );
  GTECH_XOR3 U357 ( .A(n346), .B(n348), .C(n347), .Z(n335) );
  GTECH_OAI21 U358 ( .A(n370), .B(n371), .C(n372), .Z(n347) );
  GTECH_NOT U359 ( .A(n373), .Z(n348) );
  GTECH_NAND2 U360 ( .A(I_b[3]), .B(I_a[2]), .Z(n373) );
  GTECH_NOT U361 ( .A(n344), .Z(n346) );
  GTECH_NAND2 U362 ( .A(I_b[2]), .B(I_a[3]), .Z(n344) );
  GTECH_NAND2 U363 ( .A(I_a[5]), .B(I_b[0]), .Z(n351) );
  GTECH_OAI21 U364 ( .A(n366), .B(n374), .C(n375), .Z(n353) );
  GTECH_OAI21 U365 ( .A(n364), .B(n376), .C(n365), .Z(n375) );
  GTECH_NOT U366 ( .A(n376), .Z(n366) );
  GTECH_NOT U367 ( .A(n377), .Z(n337) );
  GTECH_NAND2 U368 ( .A(I_a[4]), .B(I_b[1]), .Z(n377) );
  GTECH_NOT U369 ( .A(n378), .Z(n357) );
  GTECH_NAND3 U370 ( .A(I_a[0]), .B(n379), .C(I_b[4]), .Z(n378) );
  GTECH_XOR2 U371 ( .A(n380), .B(n379), .Z(N144) );
  GTECH_XOR2 U372 ( .A(n381), .B(n382), .Z(n379) );
  GTECH_XOR4 U373 ( .A(n365), .B(n376), .C(n363), .D(n364), .Z(n382) );
  GTECH_NOT U374 ( .A(n374), .Z(n364) );
  GTECH_NAND2 U375 ( .A(I_a[4]), .B(I_b[0]), .Z(n374) );
  GTECH_XOR3 U376 ( .A(n383), .B(n384), .C(n372), .Z(n363) );
  GTECH_NAND3 U377 ( .A(I_b[2]), .B(I_a[1]), .C(n385), .Z(n372) );
  GTECH_NOT U378 ( .A(n371), .Z(n384) );
  GTECH_NAND2 U379 ( .A(I_b[3]), .B(I_a[1]), .Z(n371) );
  GTECH_NOT U380 ( .A(n370), .Z(n383) );
  GTECH_NAND2 U381 ( .A(I_b[2]), .B(I_a[2]), .Z(n370) );
  GTECH_OAI21 U382 ( .A(n386), .B(n387), .C(n388), .Z(n376) );
  GTECH_OAI21 U383 ( .A(n389), .B(n390), .C(n391), .Z(n388) );
  GTECH_NOT U384 ( .A(n390), .Z(n386) );
  GTECH_NOT U385 ( .A(n392), .Z(n365) );
  GTECH_NAND2 U386 ( .A(I_a[3]), .B(I_b[1]), .Z(n392) );
  GTECH_OA21 U387 ( .A(n367), .B(n368), .C(n369), .Z(n381) );
  GTECH_OAI21 U388 ( .A(n393), .B(n394), .C(n395), .Z(n369) );
  GTECH_NOT U389 ( .A(n367), .Z(n394) );
  GTECH_AND2 U390 ( .A(I_b[4]), .B(I_a[0]), .Z(n380) );
  GTECH_XOR3 U391 ( .A(n395), .B(n368), .C(n367), .Z(N143) );
  GTECH_XOR2 U392 ( .A(n396), .B(n385), .Z(n367) );
  GTECH_NOT U393 ( .A(n397), .Z(n385) );
  GTECH_NAND2 U394 ( .A(I_b[3]), .B(I_a[0]), .Z(n397) );
  GTECH_NAND2 U395 ( .A(I_b[2]), .B(I_a[1]), .Z(n396) );
  GTECH_NOT U396 ( .A(n393), .Z(n368) );
  GTECH_XOR3 U397 ( .A(n389), .B(n391), .C(n390), .Z(n393) );
  GTECH_OAI21 U398 ( .A(n398), .B(n399), .C(n400), .Z(n390) );
  GTECH_NOT U399 ( .A(n401), .Z(n391) );
  GTECH_NAND2 U400 ( .A(I_b[1]), .B(I_a[2]), .Z(n401) );
  GTECH_NOT U401 ( .A(n387), .Z(n389) );
  GTECH_NAND2 U402 ( .A(I_b[0]), .B(I_a[3]), .Z(n387) );
  GTECH_NOT U403 ( .A(n402), .Z(n395) );
  GTECH_NAND3 U404 ( .A(I_a[0]), .B(n403), .C(I_b[2]), .Z(n402) );
  GTECH_XOR2 U405 ( .A(n404), .B(n403), .Z(N142) );
  GTECH_NOT U406 ( .A(n405), .Z(n403) );
  GTECH_XOR3 U407 ( .A(n406), .B(n407), .C(n400), .Z(n405) );
  GTECH_NAND3 U408 ( .A(n408), .B(I_b[0]), .C(I_a[1]), .Z(n400) );
  GTECH_NOT U409 ( .A(n398), .Z(n407) );
  GTECH_NAND2 U410 ( .A(I_a[1]), .B(I_b[1]), .Z(n398) );
  GTECH_NOT U411 ( .A(n399), .Z(n406) );
  GTECH_NAND2 U412 ( .A(I_b[0]), .B(I_a[2]), .Z(n399) );
  GTECH_AND2 U413 ( .A(I_b[2]), .B(I_a[0]), .Z(n404) );
  GTECH_XOR2 U414 ( .A(n408), .B(n409), .Z(N141) );
  GTECH_AND2 U415 ( .A(I_a[1]), .B(I_b[0]), .Z(n409) );
  GTECH_NOT U416 ( .A(n410), .Z(n408) );
  GTECH_NAND2 U417 ( .A(I_a[0]), .B(I_b[1]), .Z(n410) );
  GTECH_AND2 U418 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

