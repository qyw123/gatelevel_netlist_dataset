
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395;

  GTECH_MUX2 U141 ( .A(n280), .B(n281), .S(n282), .Z(sum[9]) );
  GTECH_AOI21 U142 ( .A(n283), .B(n284), .C(n285), .Z(n282) );
  GTECH_XOR2 U143 ( .A(b[9]), .B(a[9]), .Z(n281) );
  GTECH_OR_NOT U144 ( .A(n286), .B(n287), .Z(n280) );
  GTECH_XNOR2 U145 ( .A(n284), .B(n288), .Z(sum[8]) );
  GTECH_MUX2 U146 ( .A(n289), .B(n290), .S(n291), .Z(sum[7]) );
  GTECH_XNOR2 U147 ( .A(n292), .B(n293), .Z(n290) );
  GTECH_OA21 U148 ( .A(n294), .B(n295), .C(n296), .Z(n293) );
  GTECH_XOR2 U149 ( .A(n292), .B(n297), .Z(n289) );
  GTECH_XOR2 U150 ( .A(a[7]), .B(b[7]), .Z(n292) );
  GTECH_MUX2 U151 ( .A(n298), .B(n299), .S(n300), .Z(sum[6]) );
  GTECH_OA21 U152 ( .A(n301), .B(n291), .C(n295), .Z(n300) );
  GTECH_OA21 U153 ( .A(n302), .B(n303), .C(n304), .Z(n295) );
  GTECH_XOR2 U154 ( .A(b[6]), .B(a[6]), .Z(n299) );
  GTECH_OR_NOT U155 ( .A(n294), .B(n296), .Z(n298) );
  GTECH_NOT U156 ( .A(n305), .Z(sum[5]) );
  GTECH_MUX2 U157 ( .A(n306), .B(n307), .S(n308), .Z(n305) );
  GTECH_OR_NOT U158 ( .A(n302), .B(n304), .Z(n308) );
  GTECH_OA21 U159 ( .A(n309), .B(n291), .C(n303), .Z(n307) );
  GTECH_ADD_ABC U160 ( .A(a[4]), .B(n310), .C(b[4]), .COUT(n306) );
  GTECH_MUX2 U161 ( .A(n311), .B(n312), .S(cin), .Z(n310) );
  GTECH_OAI21 U162 ( .A(n313), .B(n314), .C(n315), .Z(n312) );
  GTECH_XOR2 U163 ( .A(n316), .B(n291), .Z(sum[4]) );
  GTECH_MUX2 U164 ( .A(n317), .B(n318), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U165 ( .A(n319), .B(n320), .Z(n318) );
  GTECH_XNOR2 U166 ( .A(n319), .B(n321), .Z(n317) );
  GTECH_OR_NOT U167 ( .A(n322), .B(n323), .Z(n321) );
  GTECH_OAI21 U168 ( .A(b[2]), .B(a[2]), .C(n324), .Z(n323) );
  GTECH_XOR2 U169 ( .A(n314), .B(b[3]), .Z(n319) );
  GTECH_MUX2 U170 ( .A(n325), .B(n326), .S(n327), .Z(sum[2]) );
  GTECH_MUX2 U171 ( .A(n328), .B(n329), .S(n324), .Z(n326) );
  GTECH_OAI21 U172 ( .A(n330), .B(n331), .C(n332), .Z(n324) );
  GTECH_MUX2 U173 ( .A(n329), .B(n328), .S(n333), .Z(n325) );
  GTECH_XNOR2 U174 ( .A(a[2]), .B(n334), .Z(n328) );
  GTECH_AO21 U175 ( .A(n334), .B(n335), .C(n322), .Z(n329) );
  GTECH_OAI21 U176 ( .A(n336), .B(n337), .C(n338), .Z(sum[1]) );
  GTECH_OAI21 U177 ( .A(n339), .B(n330), .C(n340), .Z(n338) );
  GTECH_OAI21 U178 ( .A(n341), .B(n327), .C(n331), .Z(n340) );
  GTECH_XNOR2 U179 ( .A(a[1]), .B(b[1]), .Z(n337) );
  GTECH_OA21 U180 ( .A(cin), .B(n342), .C(n343), .Z(n336) );
  GTECH_MUX2 U181 ( .A(n344), .B(n345), .S(n346), .Z(sum[15]) );
  GTECH_XNOR2 U182 ( .A(n347), .B(n348), .Z(n345) );
  GTECH_XNOR2 U183 ( .A(n347), .B(n349), .Z(n344) );
  GTECH_OA21 U184 ( .A(n350), .B(n351), .C(n352), .Z(n349) );
  GTECH_XNOR2 U185 ( .A(a[15]), .B(n353), .Z(n347) );
  GTECH_MUX2 U186 ( .A(n354), .B(n355), .S(n356), .Z(sum[14]) );
  GTECH_OA21 U187 ( .A(n357), .B(n358), .C(n351), .Z(n356) );
  GTECH_AOI21 U188 ( .A(n359), .B(n360), .C(n361), .Z(n351) );
  GTECH_XOR2 U189 ( .A(b[14]), .B(a[14]), .Z(n355) );
  GTECH_OR_NOT U190 ( .A(n350), .B(n352), .Z(n354) );
  GTECH_MUX2 U191 ( .A(n362), .B(n363), .S(n346), .Z(sum[13]) );
  GTECH_XOR2 U192 ( .A(n364), .B(n365), .Z(n363) );
  GTECH_XNOR2 U193 ( .A(n360), .B(n364), .Z(n362) );
  GTECH_OR_NOT U194 ( .A(n361), .B(n359), .Z(n364) );
  GTECH_NAND2 U195 ( .A(n366), .B(n367), .Z(sum[12]) );
  GTECH_OAI21 U196 ( .A(n365), .B(n360), .C(n346), .Z(n367) );
  GTECH_NOT U197 ( .A(n358), .Z(n346) );
  GTECH_NOT U198 ( .A(n368), .Z(n365) );
  GTECH_MUX2 U199 ( .A(n369), .B(n370), .S(n284), .Z(sum[11]) );
  GTECH_XOR2 U200 ( .A(n371), .B(n372), .Z(n370) );
  GTECH_XNOR2 U201 ( .A(n371), .B(n373), .Z(n369) );
  GTECH_OA21 U202 ( .A(n374), .B(n375), .C(n376), .Z(n373) );
  GTECH_NOT U203 ( .A(n377), .Z(n376) );
  GTECH_XOR2 U204 ( .A(a[11]), .B(b[11]), .Z(n371) );
  GTECH_MUX2 U205 ( .A(n378), .B(n379), .S(n284), .Z(sum[10]) );
  GTECH_XOR2 U206 ( .A(n380), .B(n381), .Z(n379) );
  GTECH_XNOR2 U207 ( .A(n375), .B(n380), .Z(n378) );
  GTECH_NOR2 U208 ( .A(n374), .B(n377), .Z(n380) );
  GTECH_AOI21 U209 ( .A(n287), .B(n285), .C(n286), .Z(n375) );
  GTECH_XOR2 U210 ( .A(n327), .B(n382), .Z(sum[0]) );
  GTECH_NOT U211 ( .A(cin), .Z(n327) );
  GTECH_OAI21 U212 ( .A(n383), .B(n358), .C(n366), .Z(cout) );
  GTECH_NAND3 U213 ( .A(n368), .B(n384), .C(n358), .Z(n366) );
  GTECH_NOT U214 ( .A(n360), .Z(n384) );
  GTECH_AND2 U215 ( .A(b[12]), .B(a[12]), .Z(n360) );
  GTECH_MUX2 U216 ( .A(n288), .B(n385), .S(n284), .Z(n358) );
  GTECH_MUX2 U217 ( .A(n386), .B(n387), .S(n291), .Z(n284) );
  GTECH_MUX2 U218 ( .A(n382), .B(n388), .S(cin), .Z(n291) );
  GTECH_OA21 U219 ( .A(n313), .B(n314), .C(n315), .Z(n388) );
  GTECH_OAI21 U220 ( .A(a[3]), .B(n320), .C(b[3]), .Z(n315) );
  GTECH_NOT U221 ( .A(a[3]), .Z(n314) );
  GTECH_NOT U222 ( .A(n320), .Z(n313) );
  GTECH_OR_NOT U223 ( .A(n322), .B(n389), .Z(n320) );
  GTECH_AO21 U224 ( .A(n335), .B(n334), .C(n333), .Z(n389) );
  GTECH_AOI21 U225 ( .A(n343), .B(n390), .C(n339), .Z(n333) );
  GTECH_NOT U226 ( .A(n332), .Z(n339) );
  GTECH_NAND2 U227 ( .A(b[1]), .B(a[1]), .Z(n332) );
  GTECH_NOT U228 ( .A(n330), .Z(n390) );
  GTECH_NOR2 U229 ( .A(a[1]), .B(b[1]), .Z(n330) );
  GTECH_NOT U230 ( .A(b[2]), .Z(n334) );
  GTECH_NOT U231 ( .A(a[2]), .Z(n335) );
  GTECH_AND2 U232 ( .A(b[2]), .B(a[2]), .Z(n322) );
  GTECH_NOT U233 ( .A(n311), .Z(n382) );
  GTECH_AND2 U234 ( .A(n343), .B(n331), .Z(n311) );
  GTECH_NOT U235 ( .A(n342), .Z(n331) );
  GTECH_AND2 U236 ( .A(b[0]), .B(a[0]), .Z(n342) );
  GTECH_NOT U237 ( .A(n341), .Z(n343) );
  GTECH_NOR2 U238 ( .A(a[0]), .B(b[0]), .Z(n341) );
  GTECH_NOT U239 ( .A(n316), .Z(n387) );
  GTECH_OR_NOT U240 ( .A(n309), .B(n303), .Z(n316) );
  GTECH_NAND2 U241 ( .A(b[4]), .B(a[4]), .Z(n303) );
  GTECH_OA21 U242 ( .A(a[7]), .B(n297), .C(n391), .Z(n386) );
  GTECH_AO21 U243 ( .A(n297), .B(a[7]), .C(b[7]), .Z(n391) );
  GTECH_OAI21 U244 ( .A(n301), .B(n294), .C(n296), .Z(n297) );
  GTECH_NAND2 U245 ( .A(b[6]), .B(a[6]), .Z(n296) );
  GTECH_NOR2 U246 ( .A(b[6]), .B(a[6]), .Z(n294) );
  GTECH_OA21 U247 ( .A(n302), .B(n309), .C(n304), .Z(n301) );
  GTECH_NAND2 U248 ( .A(a[5]), .B(b[5]), .Z(n304) );
  GTECH_NOR2 U249 ( .A(b[4]), .B(a[4]), .Z(n309) );
  GTECH_NOR2 U250 ( .A(a[5]), .B(b[5]), .Z(n302) );
  GTECH_AOI21 U251 ( .A(n372), .B(a[11]), .C(n392), .Z(n385) );
  GTECH_OA21 U252 ( .A(a[11]), .B(n372), .C(b[11]), .Z(n392) );
  GTECH_AO21 U253 ( .A(n381), .B(n393), .C(n377), .Z(n372) );
  GTECH_AND2 U254 ( .A(b[10]), .B(a[10]), .Z(n377) );
  GTECH_NOT U255 ( .A(n374), .Z(n393) );
  GTECH_NOR2 U256 ( .A(b[10]), .B(a[10]), .Z(n374) );
  GTECH_AO21 U257 ( .A(n283), .B(n287), .C(n286), .Z(n381) );
  GTECH_AND2 U258 ( .A(a[9]), .B(b[9]), .Z(n286) );
  GTECH_OR2 U259 ( .A(b[9]), .B(a[9]), .Z(n287) );
  GTECH_OR_NOT U260 ( .A(n285), .B(n283), .Z(n288) );
  GTECH_OR2 U261 ( .A(b[8]), .B(a[8]), .Z(n283) );
  GTECH_AND2 U262 ( .A(b[8]), .B(a[8]), .Z(n285) );
  GTECH_OA21 U263 ( .A(n348), .B(n394), .C(n395), .Z(n383) );
  GTECH_AO21 U264 ( .A(n394), .B(n348), .C(n353), .Z(n395) );
  GTECH_NOT U265 ( .A(b[15]), .Z(n353) );
  GTECH_NOT U266 ( .A(a[15]), .Z(n394) );
  GTECH_OA21 U267 ( .A(n357), .B(n350), .C(n352), .Z(n348) );
  GTECH_NAND2 U268 ( .A(b[14]), .B(a[14]), .Z(n352) );
  GTECH_NOR2 U269 ( .A(b[14]), .B(a[14]), .Z(n350) );
  GTECH_AOI21 U270 ( .A(n368), .B(n359), .C(n361), .Z(n357) );
  GTECH_AND2 U271 ( .A(a[13]), .B(b[13]), .Z(n361) );
  GTECH_OR2 U272 ( .A(a[13]), .B(b[13]), .Z(n359) );
  GTECH_OR2 U273 ( .A(b[12]), .B(a[12]), .Z(n368) );
endmodule

