
module ripple_carry_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64;

  GTECH_XNOR3 U41 ( .A(b[9]), .B(a[9]), .C(n24), .Z(sum[9]) );
  GTECH_XNOR3 U42 ( .A(b[8]), .B(a[8]), .C(n25), .Z(sum[8]) );
  GTECH_XNOR3 U43 ( .A(b[7]), .B(a[7]), .C(n26), .Z(sum[7]) );
  GTECH_XNOR3 U44 ( .A(b[6]), .B(a[6]), .C(n27), .Z(sum[6]) );
  GTECH_XNOR3 U45 ( .A(b[5]), .B(a[5]), .C(n28), .Z(sum[5]) );
  GTECH_XNOR3 U46 ( .A(b[4]), .B(a[4]), .C(n29), .Z(sum[4]) );
  GTECH_ADD_ABC U47 ( .A(b[3]), .B(a[3]), .C(n30), .S(sum[3]) );
  GTECH_XNOR3 U48 ( .A(b[2]), .B(a[2]), .C(n31), .Z(sum[2]) );
  GTECH_OAI21 U49 ( .A(a[1]), .B(n32), .C(n33), .Z(n31) );
  GTECH_ADD_ABC U50 ( .A(b[1]), .B(a[1]), .C(n32), .S(sum[1]) );
  GTECH_XNOR3 U51 ( .A(b[15]), .B(a[15]), .C(n34), .Z(sum[15]) );
  GTECH_ADD_ABC U52 ( .A(b[14]), .B(a[14]), .C(n35), .S(sum[14]) );
  GTECH_ADD_ABC U53 ( .A(b[13]), .B(a[13]), .C(n36), .S(sum[13]) );
  GTECH_ADD_ABC U54 ( .A(b[12]), .B(a[12]), .C(n37), .S(sum[12]) );
  GTECH_XNOR3 U55 ( .A(b[11]), .B(a[11]), .C(n38), .Z(sum[11]) );
  GTECH_OAI21 U56 ( .A(a[10]), .B(n39), .C(n40), .Z(n38) );
  GTECH_XNOR3 U57 ( .A(b[10]), .B(a[10]), .C(n41), .Z(sum[10]) );
  GTECH_ADD_ABC U58 ( .A(cin), .B(b[0]), .C(a[0]), .S(sum[0]) );
  GTECH_OAI21 U59 ( .A(n34), .B(n42), .C(n43), .Z(cout) );
  GTECH_OAI21 U60 ( .A(a[15]), .B(n44), .C(b[15]), .Z(n43) );
  GTECH_NOT U61 ( .A(n34), .Z(n44) );
  GTECH_NOT U62 ( .A(a[15]), .Z(n42) );
  GTECH_AOI21 U63 ( .A(n35), .B(a[14]), .C(n45), .Z(n34) );
  GTECH_OA21 U64 ( .A(a[14]), .B(n35), .C(b[14]), .Z(n45) );
  GTECH_NOT U65 ( .A(n46), .Z(n35) );
  GTECH_AOI21 U66 ( .A(n36), .B(a[13]), .C(n47), .Z(n46) );
  GTECH_OA21 U67 ( .A(a[13]), .B(n36), .C(b[13]), .Z(n47) );
  GTECH_ADD_ABC U68 ( .A(n37), .B(a[12]), .C(b[12]), .COUT(n36) );
  GTECH_ADD_ABC U69 ( .A(a[11]), .B(n48), .C(b[11]), .COUT(n37) );
  GTECH_OA21 U70 ( .A(a[10]), .B(n39), .C(n40), .Z(n48) );
  GTECH_NOT U71 ( .A(n49), .Z(n40) );
  GTECH_AOI21 U72 ( .A(n39), .B(a[10]), .C(b[10]), .Z(n49) );
  GTECH_NOT U73 ( .A(n41), .Z(n39) );
  GTECH_AOI21 U74 ( .A(n50), .B(a[9]), .C(n51), .Z(n41) );
  GTECH_OA21 U75 ( .A(a[9]), .B(n50), .C(b[9]), .Z(n51) );
  GTECH_NOT U76 ( .A(n24), .Z(n50) );
  GTECH_AOI21 U77 ( .A(n52), .B(a[8]), .C(n53), .Z(n24) );
  GTECH_OA21 U78 ( .A(a[8]), .B(n52), .C(b[8]), .Z(n53) );
  GTECH_NOT U79 ( .A(n25), .Z(n52) );
  GTECH_AOI21 U80 ( .A(n54), .B(a[7]), .C(n55), .Z(n25) );
  GTECH_OA21 U81 ( .A(a[7]), .B(n54), .C(b[7]), .Z(n55) );
  GTECH_NOT U82 ( .A(n26), .Z(n54) );
  GTECH_AOI21 U83 ( .A(n56), .B(a[6]), .C(n57), .Z(n26) );
  GTECH_OA21 U84 ( .A(a[6]), .B(n56), .C(b[6]), .Z(n57) );
  GTECH_NOT U85 ( .A(n27), .Z(n56) );
  GTECH_AOI21 U86 ( .A(n58), .B(a[5]), .C(n59), .Z(n27) );
  GTECH_OA21 U87 ( .A(a[5]), .B(n58), .C(b[5]), .Z(n59) );
  GTECH_NOT U88 ( .A(n28), .Z(n58) );
  GTECH_AOI21 U89 ( .A(n60), .B(a[4]), .C(n61), .Z(n28) );
  GTECH_OA21 U90 ( .A(a[4]), .B(n60), .C(b[4]), .Z(n61) );
  GTECH_NOT U91 ( .A(n29), .Z(n60) );
  GTECH_AOI21 U92 ( .A(n30), .B(a[3]), .C(n62), .Z(n29) );
  GTECH_OA21 U93 ( .A(a[3]), .B(n30), .C(b[3]), .Z(n62) );
  GTECH_ADD_ABC U94 ( .A(n63), .B(a[2]), .C(b[2]), .COUT(n30) );
  GTECH_OA21 U95 ( .A(a[1]), .B(n32), .C(n33), .Z(n63) );
  GTECH_NOT U96 ( .A(n64), .Z(n33) );
  GTECH_AOI21 U97 ( .A(n32), .B(a[1]), .C(b[1]), .Z(n64) );
  GTECH_ADD_ABC U98 ( .A(a[0]), .B(b[0]), .C(cin), .COUT(n32) );
endmodule

