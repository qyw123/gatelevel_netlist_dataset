
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n1, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439;

  GTECH_FD2S O_valid_reg ( .D(I_valid), .TI(n1), .TE(n1), .CP(clk), .CD(
        I_reset_n), .Q(O_valid) );
  GTECH_FD2S O_c_reg_15_ ( .D(N155), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2S O_c_reg_14_ ( .D(N154), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2S O_c_reg_13_ ( .D(N153), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2S O_c_reg_12_ ( .D(N152), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2S O_c_reg_11_ ( .D(N151), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2S O_c_reg_10_ ( .D(N150), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2S O_c_reg_9_ ( .D(N149), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[9]) );
  GTECH_FD2S O_c_reg_8_ ( .D(N148), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[8]) );
  GTECH_FD2S O_c_reg_7_ ( .D(N147), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[7]) );
  GTECH_FD2S O_c_reg_6_ ( .D(N146), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[6]) );
  GTECH_FD2S O_c_reg_5_ ( .D(N145), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[5]) );
  GTECH_FD2S O_c_reg_4_ ( .D(N144), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[4]) );
  GTECH_FD2S O_c_reg_3_ ( .D(N143), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[3]) );
  GTECH_FD2S O_c_reg_2_ ( .D(N142), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[2]) );
  GTECH_FD2S O_c_reg_1_ ( .D(N141), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[1]) );
  GTECH_FD2S O_c_reg_0_ ( .D(N140), .TI(n1), .TE(n1), .CP(clk), .CD(I_reset_n), 
        .Q(O_c[0]) );
  GTECH_ZERO U92 ( .Z(n1) );
  GTECH_NOT U93 ( .A(n100), .Z(N155) );
  GTECH_AOI222 U94 ( .A(n101), .B(n102), .C(n103), .D(n104), .E(n105), .F(n106), .Z(n100) );
  GTECH_NOT U95 ( .A(n107), .Z(n105) );
  GTECH_XOR2 U96 ( .A(n101), .B(n102), .Z(N154) );
  GTECH_NOT U97 ( .A(n108), .Z(n102) );
  GTECH_XOR2 U98 ( .A(n103), .B(n109), .Z(n108) );
  GTECH_NOT U99 ( .A(n104), .Z(n109) );
  GTECH_OAI2N2 U100 ( .A(n110), .B(n111), .C(n112), .D(n113), .Z(n104) );
  GTECH_OR_NOT U101 ( .A(n114), .B(n110), .Z(n113) );
  GTECH_XOR2 U102 ( .A(n107), .B(n115), .Z(n103) );
  GTECH_NOT U103 ( .A(n106), .Z(n115) );
  GTECH_OAI21 U104 ( .A(n116), .B(n117), .C(n118), .Z(n106) );
  GTECH_OAI21 U105 ( .A(n119), .B(n120), .C(n121), .Z(n118) );
  GTECH_NOT U106 ( .A(n120), .Z(n116) );
  GTECH_OR_NOT U107 ( .A(n122), .B(I_b[7]), .Z(n107) );
  GTECH_NOT U108 ( .A(n123), .Z(n101) );
  GTECH_OR_NOT U109 ( .A(n124), .B(n125), .Z(n123) );
  GTECH_XOR2 U110 ( .A(n126), .B(n125), .Z(N153) );
  GTECH_NOT U111 ( .A(n127), .Z(n125) );
  GTECH_XOR3 U112 ( .A(n114), .B(n110), .C(n112), .Z(n127) );
  GTECH_XOR3 U113 ( .A(n119), .B(n121), .C(n120), .Z(n112) );
  GTECH_OAI21 U114 ( .A(n128), .B(n129), .C(n130), .Z(n120) );
  GTECH_OAI21 U115 ( .A(n131), .B(n132), .C(n133), .Z(n130) );
  GTECH_NOT U116 ( .A(n132), .Z(n128) );
  GTECH_NOT U117 ( .A(n134), .Z(n121) );
  GTECH_OR_NOT U118 ( .A(n135), .B(I_b[7]), .Z(n134) );
  GTECH_NOT U119 ( .A(n117), .Z(n119) );
  GTECH_OR_NOT U120 ( .A(n136), .B(I_a[7]), .Z(n117) );
  GTECH_NOT U121 ( .A(I_b[6]), .Z(n136) );
  GTECH_ADD_ABC U122 ( .A(n137), .B(n138), .C(n139), .COUT(n110) );
  GTECH_NOT U123 ( .A(n140), .Z(n139) );
  GTECH_XOR2 U124 ( .A(n141), .B(n142), .Z(n138) );
  GTECH_AND2 U125 ( .A(I_a[7]), .B(I_b[5]), .Z(n142) );
  GTECH_NOT U126 ( .A(n111), .Z(n114) );
  GTECH_OR_NOT U127 ( .A(n141), .B(I_a[7]), .Z(n111) );
  GTECH_NOT U128 ( .A(n124), .Z(n126) );
  GTECH_OR_NOT U129 ( .A(n143), .B(n144), .Z(n124) );
  GTECH_XOR2 U130 ( .A(n143), .B(n145), .Z(N152) );
  GTECH_NOT U131 ( .A(n144), .Z(n145) );
  GTECH_XOR4 U132 ( .A(n146), .B(n141), .C(n137), .D(n140), .Z(n144) );
  GTECH_XOR3 U133 ( .A(n131), .B(n133), .C(n132), .Z(n140) );
  GTECH_OAI21 U134 ( .A(n147), .B(n148), .C(n149), .Z(n132) );
  GTECH_OAI21 U135 ( .A(n150), .B(n151), .C(n152), .Z(n149) );
  GTECH_NOT U136 ( .A(n151), .Z(n147) );
  GTECH_NOT U137 ( .A(n153), .Z(n133) );
  GTECH_OR_NOT U138 ( .A(n154), .B(I_b[7]), .Z(n153) );
  GTECH_NOT U139 ( .A(n129), .Z(n131) );
  GTECH_OR_NOT U140 ( .A(n135), .B(I_b[6]), .Z(n129) );
  GTECH_NOT U141 ( .A(I_a[6]), .Z(n135) );
  GTECH_ADD_ABC U142 ( .A(n155), .B(n156), .C(n157), .COUT(n137) );
  GTECH_NOT U143 ( .A(n158), .Z(n157) );
  GTECH_XOR3 U144 ( .A(n159), .B(n160), .C(n161), .Z(n156) );
  GTECH_OA21 U145 ( .A(n161), .B(n162), .C(n163), .Z(n141) );
  GTECH_OAI21 U146 ( .A(n159), .B(n164), .C(n160), .Z(n163) );
  GTECH_NOT U147 ( .A(n162), .Z(n159) );
  GTECH_NOT U148 ( .A(n164), .Z(n161) );
  GTECH_AND2 U149 ( .A(I_b[5]), .B(I_a[7]), .Z(n146) );
  GTECH_ADD_ABC U150 ( .A(n165), .B(n166), .C(n167), .COUT(n143) );
  GTECH_NOT U151 ( .A(n168), .Z(n167) );
  GTECH_OA22 U152 ( .A(n169), .B(n122), .C(n170), .D(n171), .Z(n166) );
  GTECH_OA21 U153 ( .A(n172), .B(n173), .C(n174), .Z(n165) );
  GTECH_XOR3 U154 ( .A(n175), .B(n168), .C(n176), .Z(N151) );
  GTECH_OA21 U155 ( .A(n172), .B(n173), .C(n174), .Z(n176) );
  GTECH_OAI21 U156 ( .A(n177), .B(n178), .C(n179), .Z(n174) );
  GTECH_XOR2 U157 ( .A(n180), .B(n155), .Z(n168) );
  GTECH_ADD_ABC U158 ( .A(n181), .B(n182), .C(n183), .COUT(n155) );
  GTECH_NOT U159 ( .A(n184), .Z(n183) );
  GTECH_XOR3 U160 ( .A(n185), .B(n186), .C(n187), .Z(n182) );
  GTECH_XOR4 U161 ( .A(n160), .B(n164), .C(n162), .D(n158), .Z(n180) );
  GTECH_XOR3 U162 ( .A(n150), .B(n152), .C(n151), .Z(n158) );
  GTECH_OAI21 U163 ( .A(n188), .B(n189), .C(n190), .Z(n151) );
  GTECH_OAI21 U164 ( .A(n191), .B(n192), .C(n193), .Z(n190) );
  GTECH_NOT U165 ( .A(n192), .Z(n188) );
  GTECH_NOT U166 ( .A(n194), .Z(n152) );
  GTECH_OR_NOT U167 ( .A(n195), .B(I_b[7]), .Z(n194) );
  GTECH_NOT U168 ( .A(n148), .Z(n150) );
  GTECH_OR_NOT U169 ( .A(n154), .B(I_b[6]), .Z(n148) );
  GTECH_NOT U170 ( .A(I_a[5]), .Z(n154) );
  GTECH_OR_NOT U171 ( .A(n196), .B(I_a[7]), .Z(n162) );
  GTECH_OAI21 U172 ( .A(n187), .B(n197), .C(n198), .Z(n164) );
  GTECH_OAI21 U173 ( .A(n185), .B(n199), .C(n186), .Z(n198) );
  GTECH_NOT U174 ( .A(n197), .Z(n185) );
  GTECH_NOT U175 ( .A(n199), .Z(n187) );
  GTECH_NOT U176 ( .A(n200), .Z(n160) );
  GTECH_OR_NOT U177 ( .A(n201), .B(I_a[6]), .Z(n200) );
  GTECH_OA22 U178 ( .A(n169), .B(n122), .C(n170), .D(n171), .Z(n175) );
  GTECH_NOT U179 ( .A(n202), .Z(n171) );
  GTECH_NOT U180 ( .A(I_a[7]), .Z(n122) );
  GTECH_XOR3 U181 ( .A(n172), .B(n177), .C(n203), .Z(N150) );
  GTECH_NOT U182 ( .A(n179), .Z(n203) );
  GTECH_XOR2 U183 ( .A(n204), .B(n181), .Z(n179) );
  GTECH_ADD_ABC U184 ( .A(n205), .B(n206), .C(n207), .COUT(n181) );
  GTECH_NOT U185 ( .A(n208), .Z(n207) );
  GTECH_XOR3 U186 ( .A(n209), .B(n210), .C(n211), .Z(n206) );
  GTECH_XOR4 U187 ( .A(n186), .B(n199), .C(n197), .D(n184), .Z(n204) );
  GTECH_XOR3 U188 ( .A(n191), .B(n193), .C(n192), .Z(n184) );
  GTECH_OAI21 U189 ( .A(n212), .B(n213), .C(n214), .Z(n192) );
  GTECH_OAI21 U190 ( .A(n215), .B(n216), .C(n217), .Z(n214) );
  GTECH_NOT U191 ( .A(n216), .Z(n212) );
  GTECH_NOT U192 ( .A(n218), .Z(n193) );
  GTECH_OR_NOT U193 ( .A(n219), .B(I_b[7]), .Z(n218) );
  GTECH_NOT U194 ( .A(n189), .Z(n191) );
  GTECH_OR_NOT U195 ( .A(n195), .B(I_b[6]), .Z(n189) );
  GTECH_OR_NOT U196 ( .A(n196), .B(I_a[6]), .Z(n197) );
  GTECH_OAI21 U197 ( .A(n211), .B(n220), .C(n221), .Z(n199) );
  GTECH_OAI21 U198 ( .A(n209), .B(n222), .C(n210), .Z(n221) );
  GTECH_NOT U199 ( .A(n220), .Z(n209) );
  GTECH_NOT U200 ( .A(n222), .Z(n211) );
  GTECH_NOT U201 ( .A(n223), .Z(n186) );
  GTECH_OR_NOT U202 ( .A(n201), .B(I_a[5]), .Z(n223) );
  GTECH_NOT U203 ( .A(I_b[5]), .Z(n201) );
  GTECH_NOT U204 ( .A(n173), .Z(n177) );
  GTECH_XOR2 U205 ( .A(n202), .B(n170), .Z(n173) );
  GTECH_AOI2N2 U206 ( .A(n224), .B(n225), .C(n226), .D(n227), .Z(n170) );
  GTECH_OR_NOT U207 ( .A(n228), .B(n226), .Z(n225) );
  GTECH_XOR2 U208 ( .A(n229), .B(n169), .Z(n202) );
  GTECH_AND2 U209 ( .A(n230), .B(n231), .Z(n169) );
  GTECH_OR_NOT U210 ( .A(n232), .B(n233), .Z(n231) );
  GTECH_OAI21 U211 ( .A(n234), .B(n233), .C(n235), .Z(n230) );
  GTECH_OR_NOT U212 ( .A(n236), .B(I_a[7]), .Z(n229) );
  GTECH_NOT U213 ( .A(n178), .Z(n172) );
  GTECH_OAI2N2 U214 ( .A(n237), .B(n238), .C(n239), .D(n240), .Z(n178) );
  GTECH_OR_NOT U215 ( .A(n241), .B(n237), .Z(n240) );
  GTECH_XOR3 U216 ( .A(n237), .B(n241), .C(n242), .Z(N149) );
  GTECH_NOT U217 ( .A(n239), .Z(n242) );
  GTECH_XOR2 U218 ( .A(n243), .B(n205), .Z(n239) );
  GTECH_ADD_ABC U219 ( .A(n244), .B(n245), .C(n246), .COUT(n205) );
  GTECH_XOR3 U220 ( .A(n247), .B(n248), .C(n249), .Z(n245) );
  GTECH_OA21 U221 ( .A(n250), .B(n251), .C(n252), .Z(n244) );
  GTECH_XOR4 U222 ( .A(n210), .B(n222), .C(n220), .D(n208), .Z(n243) );
  GTECH_XOR3 U223 ( .A(n215), .B(n217), .C(n216), .Z(n208) );
  GTECH_OAI21 U224 ( .A(n253), .B(n254), .C(n255), .Z(n216) );
  GTECH_NOT U225 ( .A(n256), .Z(n217) );
  GTECH_OR_NOT U226 ( .A(n257), .B(I_b[7]), .Z(n256) );
  GTECH_NOT U227 ( .A(n213), .Z(n215) );
  GTECH_OR_NOT U228 ( .A(n219), .B(I_b[6]), .Z(n213) );
  GTECH_OR_NOT U229 ( .A(n196), .B(I_a[5]), .Z(n220) );
  GTECH_NOT U230 ( .A(I_b[4]), .Z(n196) );
  GTECH_OAI21 U231 ( .A(n249), .B(n258), .C(n259), .Z(n222) );
  GTECH_OAI21 U232 ( .A(n247), .B(n260), .C(n248), .Z(n259) );
  GTECH_NOT U233 ( .A(n258), .Z(n247) );
  GTECH_NOT U234 ( .A(n260), .Z(n249) );
  GTECH_NOT U235 ( .A(n261), .Z(n210) );
  GTECH_OR_NOT U236 ( .A(n195), .B(I_b[5]), .Z(n261) );
  GTECH_NOT U237 ( .A(n238), .Z(n241) );
  GTECH_XOR3 U238 ( .A(n228), .B(n226), .C(n224), .Z(n238) );
  GTECH_XOR3 U239 ( .A(n234), .B(n235), .C(n233), .Z(n224) );
  GTECH_OAI21 U240 ( .A(n262), .B(n263), .C(n264), .Z(n233) );
  GTECH_OAI21 U241 ( .A(n265), .B(n266), .C(n267), .Z(n264) );
  GTECH_NOT U242 ( .A(n266), .Z(n262) );
  GTECH_NOT U243 ( .A(n268), .Z(n235) );
  GTECH_OR_NOT U244 ( .A(n236), .B(I_a[6]), .Z(n268) );
  GTECH_NOT U245 ( .A(n232), .Z(n234) );
  GTECH_OR_NOT U246 ( .A(n269), .B(I_a[7]), .Z(n232) );
  GTECH_ADD_ABC U247 ( .A(n270), .B(n271), .C(n272), .COUT(n226) );
  GTECH_XOR2 U248 ( .A(n273), .B(n274), .Z(n271) );
  GTECH_AND2 U249 ( .A(I_a[7]), .B(I_b[1]), .Z(n274) );
  GTECH_NOT U250 ( .A(n227), .Z(n228) );
  GTECH_OR_NOT U251 ( .A(n273), .B(I_a[7]), .Z(n227) );
  GTECH_ADD_ABC U252 ( .A(n275), .B(n276), .C(n277), .COUT(n237) );
  GTECH_XOR3 U253 ( .A(n270), .B(n278), .C(n272), .Z(n276) );
  GTECH_NOT U254 ( .A(n279), .Z(n272) );
  GTECH_XOR2 U255 ( .A(n275), .B(n280), .Z(N148) );
  GTECH_XOR4 U256 ( .A(n278), .B(n279), .C(n277), .D(n270), .Z(n280) );
  GTECH_ADD_ABC U257 ( .A(n281), .B(n282), .C(n283), .COUT(n270) );
  GTECH_XOR3 U258 ( .A(n284), .B(n285), .C(n286), .Z(n282) );
  GTECH_XOR2 U259 ( .A(n287), .B(n288), .Z(n277) );
  GTECH_OA21 U260 ( .A(n250), .B(n251), .C(n252), .Z(n288) );
  GTECH_OAI21 U261 ( .A(n289), .B(n290), .C(n291), .Z(n252) );
  GTECH_NOT U262 ( .A(n250), .Z(n290) );
  GTECH_XOR4 U263 ( .A(n248), .B(n260), .C(n258), .D(n246), .Z(n287) );
  GTECH_XOR3 U264 ( .A(n292), .B(n293), .C(n255), .Z(n246) );
  GTECH_NAND3 U265 ( .A(I_b[6]), .B(I_a[1]), .C(n294), .Z(n255) );
  GTECH_NOT U266 ( .A(n254), .Z(n293) );
  GTECH_OR_NOT U267 ( .A(n295), .B(I_b[7]), .Z(n254) );
  GTECH_NOT U268 ( .A(n253), .Z(n292) );
  GTECH_OR_NOT U269 ( .A(n257), .B(I_b[6]), .Z(n253) );
  GTECH_OR_NOT U270 ( .A(n195), .B(I_b[4]), .Z(n258) );
  GTECH_OAI21 U271 ( .A(n296), .B(n297), .C(n298), .Z(n260) );
  GTECH_OAI21 U272 ( .A(n299), .B(n300), .C(n301), .Z(n298) );
  GTECH_NOT U273 ( .A(n300), .Z(n296) );
  GTECH_NOT U274 ( .A(n302), .Z(n248) );
  GTECH_OR_NOT U275 ( .A(n219), .B(I_b[5]), .Z(n302) );
  GTECH_XOR3 U276 ( .A(n265), .B(n267), .C(n266), .Z(n279) );
  GTECH_OAI21 U277 ( .A(n303), .B(n304), .C(n305), .Z(n266) );
  GTECH_OAI21 U278 ( .A(n306), .B(n307), .C(n308), .Z(n305) );
  GTECH_NOT U279 ( .A(n307), .Z(n303) );
  GTECH_NOT U280 ( .A(n309), .Z(n267) );
  GTECH_OR_NOT U281 ( .A(n236), .B(I_a[5]), .Z(n309) );
  GTECH_NOT U282 ( .A(I_b[3]), .Z(n236) );
  GTECH_NOT U283 ( .A(n263), .Z(n265) );
  GTECH_OR_NOT U284 ( .A(n269), .B(I_a[6]), .Z(n263) );
  GTECH_XOR2 U285 ( .A(n310), .B(n273), .Z(n278) );
  GTECH_OA21 U286 ( .A(n286), .B(n311), .C(n312), .Z(n273) );
  GTECH_OAI21 U287 ( .A(n284), .B(n313), .C(n285), .Z(n312) );
  GTECH_NOT U288 ( .A(n313), .Z(n286) );
  GTECH_AND2 U289 ( .A(I_b[1]), .B(I_a[7]), .Z(n310) );
  GTECH_ADD_ABC U290 ( .A(n314), .B(n315), .C(n316), .COUT(n275) );
  GTECH_NOT U291 ( .A(n317), .Z(n316) );
  GTECH_XOR3 U292 ( .A(n281), .B(n318), .C(n283), .Z(n315) );
  GTECH_NOT U293 ( .A(n319), .Z(n283) );
  GTECH_NOT U294 ( .A(n320), .Z(n318) );
  GTECH_XOR2 U295 ( .A(n321), .B(n314), .Z(N147) );
  GTECH_ADD_ABC U296 ( .A(n322), .B(n323), .C(n324), .COUT(n314) );
  GTECH_XOR3 U297 ( .A(n325), .B(n326), .C(n327), .Z(n323) );
  GTECH_OA21 U298 ( .A(n328), .B(n329), .C(n330), .Z(n322) );
  GTECH_XOR4 U299 ( .A(n319), .B(n281), .C(n320), .D(n317), .Z(n321) );
  GTECH_XOR3 U300 ( .A(n291), .B(n251), .C(n250), .Z(n317) );
  GTECH_XOR2 U301 ( .A(n331), .B(n294), .Z(n250) );
  GTECH_NOT U302 ( .A(n332), .Z(n294) );
  GTECH_OR_NOT U303 ( .A(n333), .B(I_b[7]), .Z(n332) );
  GTECH_OR_NOT U304 ( .A(n295), .B(I_b[6]), .Z(n331) );
  GTECH_NOT U305 ( .A(n289), .Z(n251) );
  GTECH_XOR3 U306 ( .A(n299), .B(n301), .C(n300), .Z(n289) );
  GTECH_OAI21 U307 ( .A(n334), .B(n335), .C(n336), .Z(n300) );
  GTECH_NOT U308 ( .A(n337), .Z(n301) );
  GTECH_OR_NOT U309 ( .A(n257), .B(I_b[5]), .Z(n337) );
  GTECH_NOT U310 ( .A(n297), .Z(n299) );
  GTECH_OR_NOT U311 ( .A(n219), .B(I_b[4]), .Z(n297) );
  GTECH_NOT U312 ( .A(n338), .Z(n291) );
  GTECH_NAND3 U313 ( .A(I_a[0]), .B(n339), .C(I_b[6]), .Z(n338) );
  GTECH_NOT U314 ( .A(n340), .Z(n339) );
  GTECH_XOR3 U315 ( .A(n284), .B(n285), .C(n313), .Z(n320) );
  GTECH_OAI21 U316 ( .A(n341), .B(n342), .C(n343), .Z(n313) );
  GTECH_OAI21 U317 ( .A(n344), .B(n345), .C(n346), .Z(n343) );
  GTECH_NOT U318 ( .A(n347), .Z(n285) );
  GTECH_OR_NOT U319 ( .A(n348), .B(I_a[6]), .Z(n347) );
  GTECH_NOT U320 ( .A(n311), .Z(n284) );
  GTECH_OR_NOT U321 ( .A(n349), .B(I_a[7]), .Z(n311) );
  GTECH_ADD_ABC U322 ( .A(n325), .B(n350), .C(n327), .COUT(n281) );
  GTECH_NOT U323 ( .A(n351), .Z(n327) );
  GTECH_XOR3 U324 ( .A(n344), .B(n346), .C(n341), .Z(n350) );
  GTECH_NOT U325 ( .A(n345), .Z(n341) );
  GTECH_XOR3 U326 ( .A(n306), .B(n308), .C(n307), .Z(n319) );
  GTECH_OAI21 U327 ( .A(n352), .B(n353), .C(n354), .Z(n307) );
  GTECH_OAI21 U328 ( .A(n355), .B(n356), .C(n357), .Z(n354) );
  GTECH_NOT U329 ( .A(n356), .Z(n352) );
  GTECH_NOT U330 ( .A(n358), .Z(n308) );
  GTECH_OR_NOT U331 ( .A(n195), .B(I_b[3]), .Z(n358) );
  GTECH_NOT U332 ( .A(n304), .Z(n306) );
  GTECH_OR_NOT U333 ( .A(n269), .B(I_a[5]), .Z(n304) );
  GTECH_NOT U334 ( .A(I_b[2]), .Z(n269) );
  GTECH_XOR2 U335 ( .A(n359), .B(n360), .Z(N146) );
  GTECH_XOR4 U336 ( .A(n326), .B(n351), .C(n324), .D(n325), .Z(n360) );
  GTECH_ADD_ABC U337 ( .A(n361), .B(n362), .C(n363), .COUT(n325) );
  GTECH_NOT U338 ( .A(n364), .Z(n363) );
  GTECH_XOR3 U339 ( .A(n365), .B(n366), .C(n367), .Z(n362) );
  GTECH_XOR2 U340 ( .A(n340), .B(n368), .Z(n324) );
  GTECH_AND2 U341 ( .A(I_b[6]), .B(I_a[0]), .Z(n368) );
  GTECH_XOR3 U342 ( .A(n369), .B(n370), .C(n336), .Z(n340) );
  GTECH_NAND3 U343 ( .A(I_b[4]), .B(I_a[1]), .C(n371), .Z(n336) );
  GTECH_NOT U344 ( .A(n335), .Z(n370) );
  GTECH_OR_NOT U345 ( .A(n295), .B(I_b[5]), .Z(n335) );
  GTECH_NOT U346 ( .A(n334), .Z(n369) );
  GTECH_OR_NOT U347 ( .A(n257), .B(I_b[4]), .Z(n334) );
  GTECH_XOR3 U348 ( .A(n355), .B(n357), .C(n356), .Z(n351) );
  GTECH_OAI21 U349 ( .A(n372), .B(n373), .C(n374), .Z(n356) );
  GTECH_OAI21 U350 ( .A(n375), .B(n376), .C(n377), .Z(n374) );
  GTECH_NOT U351 ( .A(n376), .Z(n372) );
  GTECH_NOT U352 ( .A(n378), .Z(n357) );
  GTECH_OR_NOT U353 ( .A(n219), .B(I_b[3]), .Z(n378) );
  GTECH_NOT U354 ( .A(n353), .Z(n355) );
  GTECH_OR_NOT U355 ( .A(n195), .B(I_b[2]), .Z(n353) );
  GTECH_NOT U356 ( .A(I_a[4]), .Z(n195) );
  GTECH_NOT U357 ( .A(n379), .Z(n326) );
  GTECH_XOR3 U358 ( .A(n344), .B(n346), .C(n345), .Z(n379) );
  GTECH_OAI21 U359 ( .A(n367), .B(n380), .C(n381), .Z(n345) );
  GTECH_OAI21 U360 ( .A(n365), .B(n382), .C(n366), .Z(n381) );
  GTECH_NOT U361 ( .A(n380), .Z(n365) );
  GTECH_NOT U362 ( .A(n382), .Z(n367) );
  GTECH_NOT U363 ( .A(n383), .Z(n346) );
  GTECH_OR_NOT U364 ( .A(n348), .B(I_a[5]), .Z(n383) );
  GTECH_NOT U365 ( .A(n342), .Z(n344) );
  GTECH_OR_NOT U366 ( .A(n349), .B(I_a[6]), .Z(n342) );
  GTECH_OA21 U367 ( .A(n328), .B(n329), .C(n330), .Z(n359) );
  GTECH_OAI21 U368 ( .A(n384), .B(n385), .C(n386), .Z(n330) );
  GTECH_NOT U369 ( .A(n328), .Z(n385) );
  GTECH_XOR3 U370 ( .A(n386), .B(n329), .C(n328), .Z(N145) );
  GTECH_XOR2 U371 ( .A(n387), .B(n371), .Z(n328) );
  GTECH_NOT U372 ( .A(n388), .Z(n371) );
  GTECH_OR_NOT U373 ( .A(n333), .B(I_b[5]), .Z(n388) );
  GTECH_OR_NOT U374 ( .A(n295), .B(I_b[4]), .Z(n387) );
  GTECH_NOT U375 ( .A(n384), .Z(n329) );
  GTECH_XOR2 U376 ( .A(n389), .B(n361), .Z(n384) );
  GTECH_ADD_ABC U377 ( .A(n390), .B(n391), .C(n392), .COUT(n361) );
  GTECH_XOR3 U378 ( .A(n393), .B(n394), .C(n395), .Z(n391) );
  GTECH_OA21 U379 ( .A(n396), .B(n397), .C(n398), .Z(n390) );
  GTECH_XOR4 U380 ( .A(n366), .B(n382), .C(n380), .D(n364), .Z(n389) );
  GTECH_XOR3 U381 ( .A(n375), .B(n377), .C(n376), .Z(n364) );
  GTECH_OAI21 U382 ( .A(n399), .B(n400), .C(n401), .Z(n376) );
  GTECH_NOT U383 ( .A(n402), .Z(n377) );
  GTECH_OR_NOT U384 ( .A(n257), .B(I_b[3]), .Z(n402) );
  GTECH_NOT U385 ( .A(n373), .Z(n375) );
  GTECH_OR_NOT U386 ( .A(n219), .B(I_b[2]), .Z(n373) );
  GTECH_OR_NOT U387 ( .A(n349), .B(I_a[5]), .Z(n380) );
  GTECH_OAI21 U388 ( .A(n395), .B(n403), .C(n404), .Z(n382) );
  GTECH_OAI21 U389 ( .A(n393), .B(n405), .C(n394), .Z(n404) );
  GTECH_NOT U390 ( .A(n405), .Z(n395) );
  GTECH_NOT U391 ( .A(n406), .Z(n366) );
  GTECH_OR_NOT U392 ( .A(n348), .B(I_a[4]), .Z(n406) );
  GTECH_NOT U393 ( .A(n407), .Z(n386) );
  GTECH_NAND3 U394 ( .A(I_a[0]), .B(n408), .C(I_b[4]), .Z(n407) );
  GTECH_XOR2 U395 ( .A(n409), .B(n408), .Z(N144) );
  GTECH_XOR2 U396 ( .A(n410), .B(n411), .Z(n408) );
  GTECH_XOR4 U397 ( .A(n394), .B(n405), .C(n392), .D(n393), .Z(n411) );
  GTECH_NOT U398 ( .A(n403), .Z(n393) );
  GTECH_OR_NOT U399 ( .A(n349), .B(I_a[4]), .Z(n403) );
  GTECH_NOT U400 ( .A(I_b[0]), .Z(n349) );
  GTECH_XOR3 U401 ( .A(n412), .B(n413), .C(n401), .Z(n392) );
  GTECH_NAND3 U402 ( .A(I_b[2]), .B(I_a[1]), .C(n414), .Z(n401) );
  GTECH_NOT U403 ( .A(n400), .Z(n413) );
  GTECH_OR_NOT U404 ( .A(n295), .B(I_b[3]), .Z(n400) );
  GTECH_NOT U405 ( .A(n399), .Z(n412) );
  GTECH_OR_NOT U406 ( .A(n257), .B(I_b[2]), .Z(n399) );
  GTECH_OAI21 U407 ( .A(n415), .B(n416), .C(n417), .Z(n405) );
  GTECH_OAI21 U408 ( .A(n418), .B(n419), .C(n420), .Z(n417) );
  GTECH_NOT U409 ( .A(n419), .Z(n415) );
  GTECH_NOT U410 ( .A(n421), .Z(n394) );
  GTECH_OR_NOT U411 ( .A(n348), .B(I_a[3]), .Z(n421) );
  GTECH_OA21 U412 ( .A(n396), .B(n397), .C(n398), .Z(n410) );
  GTECH_OAI21 U413 ( .A(n422), .B(n423), .C(n424), .Z(n398) );
  GTECH_NOT U414 ( .A(n396), .Z(n423) );
  GTECH_AND2 U415 ( .A(I_b[4]), .B(I_a[0]), .Z(n409) );
  GTECH_XOR3 U416 ( .A(n424), .B(n397), .C(n396), .Z(N143) );
  GTECH_XOR2 U417 ( .A(n425), .B(n414), .Z(n396) );
  GTECH_NOT U418 ( .A(n426), .Z(n414) );
  GTECH_OR_NOT U419 ( .A(n333), .B(I_b[3]), .Z(n426) );
  GTECH_NOT U420 ( .A(I_a[0]), .Z(n333) );
  GTECH_OR_NOT U421 ( .A(n295), .B(I_b[2]), .Z(n425) );
  GTECH_NOT U422 ( .A(I_a[1]), .Z(n295) );
  GTECH_NOT U423 ( .A(n422), .Z(n397) );
  GTECH_XOR3 U424 ( .A(n418), .B(n420), .C(n419), .Z(n422) );
  GTECH_OAI21 U425 ( .A(n427), .B(n428), .C(n429), .Z(n419) );
  GTECH_NOT U426 ( .A(n430), .Z(n420) );
  GTECH_OR_NOT U427 ( .A(n257), .B(I_b[1]), .Z(n430) );
  GTECH_NOT U428 ( .A(n416), .Z(n418) );
  GTECH_OR_NOT U429 ( .A(n219), .B(I_b[0]), .Z(n416) );
  GTECH_NOT U430 ( .A(I_a[3]), .Z(n219) );
  GTECH_NOT U431 ( .A(n431), .Z(n424) );
  GTECH_NAND3 U432 ( .A(I_a[0]), .B(n432), .C(I_b[2]), .Z(n431) );
  GTECH_XOR2 U433 ( .A(n433), .B(n432), .Z(N142) );
  GTECH_NOT U434 ( .A(n434), .Z(n432) );
  GTECH_XOR3 U435 ( .A(n435), .B(n436), .C(n429), .Z(n434) );
  GTECH_NAND3 U436 ( .A(n437), .B(I_b[0]), .C(I_a[1]), .Z(n429) );
  GTECH_NOT U437 ( .A(n427), .Z(n436) );
  GTECH_OR_NOT U438 ( .A(n348), .B(I_a[1]), .Z(n427) );
  GTECH_NOT U439 ( .A(n428), .Z(n435) );
  GTECH_OR_NOT U440 ( .A(n257), .B(I_b[0]), .Z(n428) );
  GTECH_NOT U441 ( .A(I_a[2]), .Z(n257) );
  GTECH_AND2 U442 ( .A(I_b[2]), .B(I_a[0]), .Z(n433) );
  GTECH_XOR2 U443 ( .A(n437), .B(n438), .Z(N141) );
  GTECH_AND2 U444 ( .A(I_a[1]), .B(I_b[0]), .Z(n438) );
  GTECH_NOT U445 ( .A(n439), .Z(n437) );
  GTECH_OR_NOT U446 ( .A(n348), .B(I_a[0]), .Z(n439) );
  GTECH_NOT U447 ( .A(I_b[1]), .Z(n348) );
  GTECH_AND2 U448 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

