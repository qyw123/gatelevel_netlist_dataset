
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NAND2 U83 ( .A(n93), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI22 U86 ( .A(n98), .B(n99), .C(n100), .D(n101), .Z(n89) );
  GTECH_AND2 U87 ( .A(n98), .B(n99), .Z(n100) );
  GTECH_NOT U88 ( .A(n102), .Z(n98) );
  GTECH_NAND2 U89 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n103), .Z(n84) );
  GTECH_NAND2 U91 ( .A(n104), .B(n105), .Z(n103) );
  GTECH_XOR2 U92 ( .A(n105), .B(n104), .Z(N153) );
  GTECH_NOT U93 ( .A(n106), .Z(n104) );
  GTECH_XOR3 U94 ( .A(n107), .B(n93), .C(n95), .Z(n106) );
  GTECH_XOR3 U95 ( .A(n108), .B(n109), .C(n102), .Z(n95) );
  GTECH_OAI22 U96 ( .A(n110), .B(n111), .C(n112), .D(n113), .Z(n102) );
  GTECH_AND2 U97 ( .A(n110), .B(n111), .Z(n112) );
  GTECH_NOT U98 ( .A(n114), .Z(n110) );
  GTECH_NOT U99 ( .A(n101), .Z(n109) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n101) );
  GTECH_NOT U101 ( .A(n99), .Z(n108) );
  GTECH_NAND2 U102 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U103 ( .A(n115), .B(n116), .C(n117), .COUT(n93) );
  GTECH_NOT U104 ( .A(n118), .Z(n117) );
  GTECH_XOR2 U105 ( .A(n119), .B(n120), .Z(n116) );
  GTECH_AND2 U106 ( .A(I_a[7]), .B(I_b[5]), .Z(n120) );
  GTECH_NOT U107 ( .A(n94), .Z(n107) );
  GTECH_NAND2 U108 ( .A(I_a[7]), .B(n121), .Z(n94) );
  GTECH_NOT U109 ( .A(n122), .Z(n105) );
  GTECH_NAND2 U110 ( .A(n123), .B(n124), .Z(n122) );
  GTECH_NOT U111 ( .A(n125), .Z(n124) );
  GTECH_XOR2 U112 ( .A(n125), .B(n126), .Z(N152) );
  GTECH_NOT U113 ( .A(n123), .Z(n126) );
  GTECH_XOR4 U114 ( .A(n127), .B(n119), .C(n115), .D(n118), .Z(n123) );
  GTECH_XOR3 U115 ( .A(n128), .B(n129), .C(n114), .Z(n118) );
  GTECH_OAI22 U116 ( .A(n130), .B(n131), .C(n132), .D(n133), .Z(n114) );
  GTECH_AND2 U117 ( .A(n130), .B(n131), .Z(n132) );
  GTECH_NOT U118 ( .A(n134), .Z(n130) );
  GTECH_NOT U119 ( .A(n113), .Z(n129) );
  GTECH_NAND2 U120 ( .A(I_b[7]), .B(I_a[5]), .Z(n113) );
  GTECH_NOT U121 ( .A(n111), .Z(n128) );
  GTECH_NAND2 U122 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_ADD_ABC U123 ( .A(n135), .B(n136), .C(n137), .COUT(n115) );
  GTECH_NOT U124 ( .A(n138), .Z(n137) );
  GTECH_XOR3 U125 ( .A(n139), .B(n140), .C(n141), .Z(n136) );
  GTECH_NOT U126 ( .A(n142), .Z(n139) );
  GTECH_NOT U127 ( .A(n121), .Z(n119) );
  GTECH_OAI22 U128 ( .A(n141), .B(n142), .C(n143), .D(n144), .Z(n121) );
  GTECH_AND2 U129 ( .A(n141), .B(n142), .Z(n143) );
  GTECH_NOT U130 ( .A(n145), .Z(n141) );
  GTECH_AND2 U131 ( .A(I_a[7]), .B(I_b[5]), .Z(n127) );
  GTECH_ADD_ABC U132 ( .A(n146), .B(n147), .C(n148), .COUT(n125) );
  GTECH_NOT U133 ( .A(n149), .Z(n148) );
  GTECH_OA22 U134 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n147) );
  GTECH_OA22 U135 ( .A(n154), .B(n155), .C(n156), .D(n157), .Z(n146) );
  GTECH_XOR3 U136 ( .A(n158), .B(n149), .C(n159), .Z(N151) );
  GTECH_OA22 U137 ( .A(n154), .B(n155), .C(n156), .D(n157), .Z(n159) );
  GTECH_AND2 U138 ( .A(n156), .B(n157), .Z(n154) );
  GTECH_XOR2 U139 ( .A(n160), .B(n135), .Z(n149) );
  GTECH_ADD_ABC U140 ( .A(n161), .B(n162), .C(n163), .COUT(n135) );
  GTECH_NOT U141 ( .A(n164), .Z(n163) );
  GTECH_XOR3 U142 ( .A(n165), .B(n166), .C(n167), .Z(n162) );
  GTECH_XOR4 U143 ( .A(n140), .B(n145), .C(n142), .D(n138), .Z(n160) );
  GTECH_XOR3 U144 ( .A(n168), .B(n169), .C(n134), .Z(n138) );
  GTECH_OAI22 U145 ( .A(n170), .B(n171), .C(n172), .D(n173), .Z(n134) );
  GTECH_AND2 U146 ( .A(n170), .B(n171), .Z(n172) );
  GTECH_NOT U147 ( .A(n174), .Z(n170) );
  GTECH_NOT U148 ( .A(n133), .Z(n169) );
  GTECH_NAND2 U149 ( .A(I_b[7]), .B(I_a[4]), .Z(n133) );
  GTECH_NOT U150 ( .A(n131), .Z(n168) );
  GTECH_NAND2 U151 ( .A(I_b[6]), .B(I_a[5]), .Z(n131) );
  GTECH_NAND2 U152 ( .A(I_a[7]), .B(I_b[4]), .Z(n142) );
  GTECH_OAI22 U153 ( .A(n167), .B(n175), .C(n176), .D(n177), .Z(n145) );
  GTECH_AND2 U154 ( .A(n167), .B(n175), .Z(n176) );
  GTECH_NOT U155 ( .A(n178), .Z(n167) );
  GTECH_NOT U156 ( .A(n144), .Z(n140) );
  GTECH_NAND2 U157 ( .A(I_a[6]), .B(I_b[5]), .Z(n144) );
  GTECH_OA22 U158 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n158) );
  GTECH_NOT U159 ( .A(n179), .Z(n153) );
  GTECH_NOT U160 ( .A(I_a[7]), .Z(n151) );
  GTECH_XOR3 U161 ( .A(n156), .B(n180), .C(n155), .Z(N150) );
  GTECH_XOR2 U162 ( .A(n161), .B(n181), .Z(n155) );
  GTECH_XOR4 U163 ( .A(n166), .B(n178), .C(n164), .D(n165), .Z(n181) );
  GTECH_NOT U164 ( .A(n175), .Z(n165) );
  GTECH_NAND2 U165 ( .A(I_a[6]), .B(I_b[4]), .Z(n175) );
  GTECH_XOR3 U166 ( .A(n182), .B(n183), .C(n174), .Z(n164) );
  GTECH_OAI22 U167 ( .A(n184), .B(n185), .C(n186), .D(n187), .Z(n174) );
  GTECH_AND2 U168 ( .A(n184), .B(n185), .Z(n186) );
  GTECH_NOT U169 ( .A(n188), .Z(n184) );
  GTECH_NOT U170 ( .A(n173), .Z(n183) );
  GTECH_NAND2 U171 ( .A(I_b[7]), .B(I_a[3]), .Z(n173) );
  GTECH_NOT U172 ( .A(n171), .Z(n182) );
  GTECH_NAND2 U173 ( .A(I_b[6]), .B(I_a[4]), .Z(n171) );
  GTECH_OAI22 U174 ( .A(n189), .B(n190), .C(n191), .D(n192), .Z(n178) );
  GTECH_AND2 U175 ( .A(n189), .B(n190), .Z(n191) );
  GTECH_NOT U176 ( .A(n177), .Z(n166) );
  GTECH_NAND2 U177 ( .A(I_a[5]), .B(I_b[5]), .Z(n177) );
  GTECH_ADD_ABC U178 ( .A(n193), .B(n194), .C(n195), .COUT(n161) );
  GTECH_NOT U179 ( .A(n196), .Z(n195) );
  GTECH_XOR3 U180 ( .A(n197), .B(n198), .C(n189), .Z(n194) );
  GTECH_NOT U181 ( .A(n199), .Z(n189) );
  GTECH_NOT U182 ( .A(n157), .Z(n180) );
  GTECH_XOR2 U183 ( .A(n179), .B(n152), .Z(n157) );
  GTECH_AOI2N2 U184 ( .A(n200), .B(n201), .C(n202), .D(n203), .Z(n152) );
  GTECH_NAND2 U185 ( .A(n202), .B(n203), .Z(n201) );
  GTECH_XOR2 U186 ( .A(n204), .B(n150), .Z(n179) );
  GTECH_OA22 U187 ( .A(n205), .B(n206), .C(n207), .D(n208), .Z(n150) );
  GTECH_AND2 U188 ( .A(n207), .B(n208), .Z(n205) );
  GTECH_NOT U189 ( .A(n209), .Z(n207) );
  GTECH_NAND2 U190 ( .A(I_a[7]), .B(I_b[3]), .Z(n204) );
  GTECH_OA22 U191 ( .A(n210), .B(n211), .C(n212), .D(n213), .Z(n156) );
  GTECH_AND2 U192 ( .A(n212), .B(n213), .Z(n210) );
  GTECH_XOR3 U193 ( .A(n212), .B(n214), .C(n211), .Z(N149) );
  GTECH_XOR2 U194 ( .A(n193), .B(n215), .Z(n211) );
  GTECH_XOR4 U195 ( .A(n198), .B(n199), .C(n196), .D(n197), .Z(n215) );
  GTECH_NOT U196 ( .A(n190), .Z(n197) );
  GTECH_NAND2 U197 ( .A(I_a[5]), .B(I_b[4]), .Z(n190) );
  GTECH_XOR3 U198 ( .A(n216), .B(n217), .C(n188), .Z(n196) );
  GTECH_AO21 U199 ( .A(n218), .B(n219), .C(n220), .Z(n188) );
  GTECH_NOT U200 ( .A(n221), .Z(n220) );
  GTECH_NOT U201 ( .A(n187), .Z(n217) );
  GTECH_NAND2 U202 ( .A(I_b[7]), .B(I_a[2]), .Z(n187) );
  GTECH_NOT U203 ( .A(n185), .Z(n216) );
  GTECH_NAND2 U204 ( .A(I_b[6]), .B(I_a[3]), .Z(n185) );
  GTECH_OAI22 U205 ( .A(n222), .B(n223), .C(n224), .D(n225), .Z(n199) );
  GTECH_AND2 U206 ( .A(n222), .B(n223), .Z(n224) );
  GTECH_NOT U207 ( .A(n192), .Z(n198) );
  GTECH_NAND2 U208 ( .A(I_b[5]), .B(I_a[4]), .Z(n192) );
  GTECH_ADD_ABC U209 ( .A(n226), .B(n227), .C(n228), .COUT(n193) );
  GTECH_XOR3 U210 ( .A(n229), .B(n230), .C(n222), .Z(n227) );
  GTECH_NOT U211 ( .A(n231), .Z(n222) );
  GTECH_NOT U212 ( .A(n223), .Z(n229) );
  GTECH_OA22 U213 ( .A(n232), .B(n233), .C(n234), .D(n235), .Z(n226) );
  GTECH_NOT U214 ( .A(n213), .Z(n214) );
  GTECH_XOR3 U215 ( .A(n236), .B(n202), .C(n200), .Z(n213) );
  GTECH_XOR3 U216 ( .A(n237), .B(n238), .C(n209), .Z(n200) );
  GTECH_OAI22 U217 ( .A(n239), .B(n240), .C(n241), .D(n242), .Z(n209) );
  GTECH_AND2 U218 ( .A(n239), .B(n240), .Z(n241) );
  GTECH_NOT U219 ( .A(n243), .Z(n239) );
  GTECH_NOT U220 ( .A(n206), .Z(n238) );
  GTECH_NAND2 U221 ( .A(I_a[6]), .B(I_b[3]), .Z(n206) );
  GTECH_NOT U222 ( .A(n208), .Z(n237) );
  GTECH_NAND2 U223 ( .A(I_a[7]), .B(I_b[2]), .Z(n208) );
  GTECH_ADD_ABC U224 ( .A(n244), .B(n245), .C(n246), .COUT(n202) );
  GTECH_XOR2 U225 ( .A(n247), .B(n248), .Z(n245) );
  GTECH_AND2 U226 ( .A(I_a[7]), .B(I_b[1]), .Z(n248) );
  GTECH_NOT U227 ( .A(n203), .Z(n236) );
  GTECH_NAND2 U228 ( .A(I_a[7]), .B(n249), .Z(n203) );
  GTECH_ADD_ABC U229 ( .A(n250), .B(n251), .C(n252), .COUT(n212) );
  GTECH_XOR3 U230 ( .A(n244), .B(n253), .C(n246), .Z(n251) );
  GTECH_NOT U231 ( .A(n254), .Z(n246) );
  GTECH_XOR2 U232 ( .A(n250), .B(n255), .Z(N148) );
  GTECH_XOR4 U233 ( .A(n253), .B(n254), .C(n252), .D(n244), .Z(n255) );
  GTECH_ADD_ABC U234 ( .A(n256), .B(n257), .C(n258), .COUT(n244) );
  GTECH_XOR3 U235 ( .A(n259), .B(n260), .C(n261), .Z(n257) );
  GTECH_XOR2 U236 ( .A(n262), .B(n263), .Z(n252) );
  GTECH_OA22 U237 ( .A(n232), .B(n233), .C(n234), .D(n235), .Z(n263) );
  GTECH_AND2 U238 ( .A(n234), .B(n235), .Z(n232) );
  GTECH_XOR4 U239 ( .A(n230), .B(n231), .C(n223), .D(n228), .Z(n262) );
  GTECH_XOR3 U240 ( .A(n219), .B(n218), .C(n221), .Z(n228) );
  GTECH_NAND3 U241 ( .A(I_b[6]), .B(I_a[1]), .C(n264), .Z(n221) );
  GTECH_NOT U242 ( .A(n265), .Z(n218) );
  GTECH_NAND2 U243 ( .A(I_b[7]), .B(I_a[1]), .Z(n265) );
  GTECH_NOT U244 ( .A(n266), .Z(n219) );
  GTECH_NAND2 U245 ( .A(I_b[6]), .B(I_a[2]), .Z(n266) );
  GTECH_NAND2 U246 ( .A(I_b[4]), .B(I_a[4]), .Z(n223) );
  GTECH_OAI22 U247 ( .A(n267), .B(n268), .C(n269), .D(n270), .Z(n231) );
  GTECH_AND2 U248 ( .A(n267), .B(n268), .Z(n269) );
  GTECH_NOT U249 ( .A(n271), .Z(n267) );
  GTECH_NOT U250 ( .A(n225), .Z(n230) );
  GTECH_NAND2 U251 ( .A(I_b[5]), .B(I_a[3]), .Z(n225) );
  GTECH_XOR3 U252 ( .A(n272), .B(n273), .C(n243), .Z(n254) );
  GTECH_OAI22 U253 ( .A(n274), .B(n275), .C(n276), .D(n277), .Z(n243) );
  GTECH_AND2 U254 ( .A(n274), .B(n275), .Z(n276) );
  GTECH_NOT U255 ( .A(n278), .Z(n274) );
  GTECH_NOT U256 ( .A(n242), .Z(n273) );
  GTECH_NAND2 U257 ( .A(I_a[5]), .B(I_b[3]), .Z(n242) );
  GTECH_NOT U258 ( .A(n240), .Z(n272) );
  GTECH_NAND2 U259 ( .A(I_a[6]), .B(I_b[2]), .Z(n240) );
  GTECH_XOR2 U260 ( .A(n279), .B(n247), .Z(n253) );
  GTECH_NOT U261 ( .A(n249), .Z(n247) );
  GTECH_OAI22 U262 ( .A(n261), .B(n280), .C(n281), .D(n282), .Z(n249) );
  GTECH_AND2 U263 ( .A(n261), .B(n280), .Z(n281) );
  GTECH_NOT U264 ( .A(n283), .Z(n261) );
  GTECH_AND2 U265 ( .A(I_a[7]), .B(I_b[1]), .Z(n279) );
  GTECH_ADD_ABC U266 ( .A(n284), .B(n285), .C(n286), .COUT(n250) );
  GTECH_NOT U267 ( .A(n287), .Z(n286) );
  GTECH_XOR3 U268 ( .A(n256), .B(n288), .C(n258), .Z(n285) );
  GTECH_NOT U269 ( .A(n289), .Z(n258) );
  GTECH_NOT U270 ( .A(n290), .Z(n288) );
  GTECH_XOR2 U271 ( .A(n291), .B(n284), .Z(N147) );
  GTECH_ADD_ABC U272 ( .A(n292), .B(n293), .C(n294), .COUT(n284) );
  GTECH_XOR3 U273 ( .A(n295), .B(n296), .C(n297), .Z(n293) );
  GTECH_OA22 U274 ( .A(n298), .B(n299), .C(n300), .D(n301), .Z(n292) );
  GTECH_XOR4 U275 ( .A(n289), .B(n256), .C(n290), .D(n287), .Z(n291) );
  GTECH_XOR3 U276 ( .A(n302), .B(n235), .C(n234), .Z(n287) );
  GTECH_XOR2 U277 ( .A(n303), .B(n264), .Z(n234) );
  GTECH_NOT U278 ( .A(n304), .Z(n264) );
  GTECH_NAND2 U279 ( .A(I_b[7]), .B(I_a[0]), .Z(n304) );
  GTECH_NAND2 U280 ( .A(I_b[6]), .B(I_a[1]), .Z(n303) );
  GTECH_NOT U281 ( .A(n305), .Z(n235) );
  GTECH_XOR3 U282 ( .A(n306), .B(n307), .C(n271), .Z(n305) );
  GTECH_AO21 U283 ( .A(n308), .B(n309), .C(n310), .Z(n271) );
  GTECH_NOT U284 ( .A(n311), .Z(n310) );
  GTECH_NOT U285 ( .A(n270), .Z(n307) );
  GTECH_NAND2 U286 ( .A(I_b[5]), .B(I_a[2]), .Z(n270) );
  GTECH_NOT U287 ( .A(n268), .Z(n306) );
  GTECH_NAND2 U288 ( .A(I_b[4]), .B(I_a[3]), .Z(n268) );
  GTECH_NOT U289 ( .A(n233), .Z(n302) );
  GTECH_NAND3 U290 ( .A(I_a[0]), .B(n312), .C(I_b[6]), .Z(n233) );
  GTECH_NOT U291 ( .A(n313), .Z(n312) );
  GTECH_XOR3 U292 ( .A(n259), .B(n260), .C(n283), .Z(n290) );
  GTECH_OAI22 U293 ( .A(n314), .B(n315), .C(n316), .D(n317), .Z(n283) );
  GTECH_AND2 U294 ( .A(n314), .B(n315), .Z(n316) );
  GTECH_NOT U295 ( .A(n282), .Z(n260) );
  GTECH_NAND2 U296 ( .A(I_a[6]), .B(I_b[1]), .Z(n282) );
  GTECH_NOT U297 ( .A(n280), .Z(n259) );
  GTECH_NAND2 U298 ( .A(I_a[7]), .B(I_b[0]), .Z(n280) );
  GTECH_ADD_ABC U299 ( .A(n295), .B(n318), .C(n297), .COUT(n256) );
  GTECH_NOT U300 ( .A(n319), .Z(n297) );
  GTECH_XOR3 U301 ( .A(n320), .B(n321), .C(n314), .Z(n318) );
  GTECH_NOT U302 ( .A(n322), .Z(n314) );
  GTECH_XOR3 U303 ( .A(n323), .B(n324), .C(n278), .Z(n289) );
  GTECH_OAI22 U304 ( .A(n325), .B(n326), .C(n327), .D(n328), .Z(n278) );
  GTECH_AND2 U305 ( .A(n325), .B(n326), .Z(n327) );
  GTECH_NOT U306 ( .A(n329), .Z(n325) );
  GTECH_NOT U307 ( .A(n277), .Z(n324) );
  GTECH_NAND2 U308 ( .A(I_b[3]), .B(I_a[4]), .Z(n277) );
  GTECH_NOT U309 ( .A(n275), .Z(n323) );
  GTECH_NAND2 U310 ( .A(I_a[5]), .B(I_b[2]), .Z(n275) );
  GTECH_XOR2 U311 ( .A(n330), .B(n331), .Z(N146) );
  GTECH_XOR4 U312 ( .A(n296), .B(n319), .C(n294), .D(n295), .Z(n331) );
  GTECH_ADD_ABC U313 ( .A(n332), .B(n333), .C(n334), .COUT(n295) );
  GTECH_NOT U314 ( .A(n335), .Z(n334) );
  GTECH_XOR3 U315 ( .A(n336), .B(n337), .C(n338), .Z(n333) );
  GTECH_XOR2 U316 ( .A(n313), .B(n339), .Z(n294) );
  GTECH_AND2 U317 ( .A(I_b[6]), .B(I_a[0]), .Z(n339) );
  GTECH_XOR3 U318 ( .A(n309), .B(n308), .C(n311), .Z(n313) );
  GTECH_NAND3 U319 ( .A(I_b[4]), .B(I_a[1]), .C(n340), .Z(n311) );
  GTECH_NOT U320 ( .A(n341), .Z(n308) );
  GTECH_NAND2 U321 ( .A(I_b[5]), .B(I_a[1]), .Z(n341) );
  GTECH_NOT U322 ( .A(n342), .Z(n309) );
  GTECH_NAND2 U323 ( .A(I_b[4]), .B(I_a[2]), .Z(n342) );
  GTECH_XOR3 U324 ( .A(n343), .B(n344), .C(n329), .Z(n319) );
  GTECH_OAI22 U325 ( .A(n345), .B(n346), .C(n347), .D(n348), .Z(n329) );
  GTECH_AND2 U326 ( .A(n345), .B(n346), .Z(n347) );
  GTECH_NOT U327 ( .A(n349), .Z(n345) );
  GTECH_NOT U328 ( .A(n328), .Z(n344) );
  GTECH_NAND2 U329 ( .A(I_b[3]), .B(I_a[3]), .Z(n328) );
  GTECH_NOT U330 ( .A(n326), .Z(n343) );
  GTECH_NAND2 U331 ( .A(I_b[2]), .B(I_a[4]), .Z(n326) );
  GTECH_NOT U332 ( .A(n350), .Z(n296) );
  GTECH_XOR3 U333 ( .A(n320), .B(n321), .C(n322), .Z(n350) );
  GTECH_OAI22 U334 ( .A(n338), .B(n351), .C(n352), .D(n353), .Z(n322) );
  GTECH_AND2 U335 ( .A(n338), .B(n351), .Z(n352) );
  GTECH_NOT U336 ( .A(n354), .Z(n338) );
  GTECH_NOT U337 ( .A(n317), .Z(n321) );
  GTECH_NAND2 U338 ( .A(I_a[5]), .B(I_b[1]), .Z(n317) );
  GTECH_NOT U339 ( .A(n315), .Z(n320) );
  GTECH_NAND2 U340 ( .A(I_a[6]), .B(I_b[0]), .Z(n315) );
  GTECH_OA22 U341 ( .A(n298), .B(n299), .C(n300), .D(n301), .Z(n330) );
  GTECH_AND2 U342 ( .A(n300), .B(n301), .Z(n298) );
  GTECH_XOR3 U343 ( .A(n355), .B(n301), .C(n300), .Z(N145) );
  GTECH_XOR2 U344 ( .A(n356), .B(n340), .Z(n300) );
  GTECH_NOT U345 ( .A(n357), .Z(n340) );
  GTECH_NAND2 U346 ( .A(I_b[5]), .B(I_a[0]), .Z(n357) );
  GTECH_NAND2 U347 ( .A(I_b[4]), .B(I_a[1]), .Z(n356) );
  GTECH_XOR2 U348 ( .A(n332), .B(n358), .Z(n301) );
  GTECH_XOR4 U349 ( .A(n337), .B(n354), .C(n335), .D(n336), .Z(n358) );
  GTECH_NOT U350 ( .A(n351), .Z(n336) );
  GTECH_NAND2 U351 ( .A(I_a[5]), .B(I_b[0]), .Z(n351) );
  GTECH_XOR3 U352 ( .A(n359), .B(n360), .C(n349), .Z(n335) );
  GTECH_AO21 U353 ( .A(n361), .B(n362), .C(n363), .Z(n349) );
  GTECH_NOT U354 ( .A(n364), .Z(n363) );
  GTECH_NOT U355 ( .A(n348), .Z(n360) );
  GTECH_NAND2 U356 ( .A(I_b[3]), .B(I_a[2]), .Z(n348) );
  GTECH_NOT U357 ( .A(n346), .Z(n359) );
  GTECH_NAND2 U358 ( .A(I_b[2]), .B(I_a[3]), .Z(n346) );
  GTECH_OAI22 U359 ( .A(n365), .B(n366), .C(n367), .D(n368), .Z(n354) );
  GTECH_AND2 U360 ( .A(n365), .B(n366), .Z(n367) );
  GTECH_NOT U361 ( .A(n353), .Z(n337) );
  GTECH_NAND2 U362 ( .A(I_a[4]), .B(I_b[1]), .Z(n353) );
  GTECH_ADD_ABC U363 ( .A(n369), .B(n370), .C(n371), .COUT(n332) );
  GTECH_XOR3 U364 ( .A(n372), .B(n373), .C(n365), .Z(n370) );
  GTECH_NOT U365 ( .A(n374), .Z(n365) );
  GTECH_OA22 U366 ( .A(n375), .B(n376), .C(n377), .D(n378), .Z(n369) );
  GTECH_NOT U367 ( .A(n299), .Z(n355) );
  GTECH_NAND3 U368 ( .A(I_a[0]), .B(n379), .C(I_b[4]), .Z(n299) );
  GTECH_XOR2 U369 ( .A(n380), .B(n379), .Z(N144) );
  GTECH_XOR2 U370 ( .A(n381), .B(n382), .Z(n379) );
  GTECH_XOR4 U371 ( .A(n373), .B(n374), .C(n371), .D(n372), .Z(n382) );
  GTECH_NOT U372 ( .A(n366), .Z(n372) );
  GTECH_NAND2 U373 ( .A(I_a[4]), .B(I_b[0]), .Z(n366) );
  GTECH_XOR3 U374 ( .A(n362), .B(n361), .C(n364), .Z(n371) );
  GTECH_NAND3 U375 ( .A(I_b[2]), .B(I_a[1]), .C(n383), .Z(n364) );
  GTECH_NOT U376 ( .A(n384), .Z(n361) );
  GTECH_NAND2 U377 ( .A(I_b[3]), .B(I_a[1]), .Z(n384) );
  GTECH_NOT U378 ( .A(n385), .Z(n362) );
  GTECH_NAND2 U379 ( .A(I_b[2]), .B(I_a[2]), .Z(n385) );
  GTECH_OAI22 U380 ( .A(n386), .B(n387), .C(n388), .D(n389), .Z(n374) );
  GTECH_AND2 U381 ( .A(n386), .B(n387), .Z(n388) );
  GTECH_NOT U382 ( .A(n390), .Z(n386) );
  GTECH_NOT U383 ( .A(n368), .Z(n373) );
  GTECH_NAND2 U384 ( .A(I_a[3]), .B(I_b[1]), .Z(n368) );
  GTECH_OA22 U385 ( .A(n375), .B(n376), .C(n377), .D(n378), .Z(n381) );
  GTECH_AND2 U386 ( .A(n377), .B(n378), .Z(n375) );
  GTECH_AND2 U387 ( .A(I_b[4]), .B(I_a[0]), .Z(n380) );
  GTECH_XOR3 U388 ( .A(n391), .B(n378), .C(n377), .Z(N143) );
  GTECH_XOR2 U389 ( .A(n392), .B(n383), .Z(n377) );
  GTECH_NOT U390 ( .A(n393), .Z(n383) );
  GTECH_NAND2 U391 ( .A(I_b[3]), .B(I_a[0]), .Z(n393) );
  GTECH_NAND2 U392 ( .A(I_b[2]), .B(I_a[1]), .Z(n392) );
  GTECH_NOT U393 ( .A(n394), .Z(n378) );
  GTECH_XOR3 U394 ( .A(n395), .B(n396), .C(n390), .Z(n394) );
  GTECH_AO21 U395 ( .A(n397), .B(n398), .C(n399), .Z(n390) );
  GTECH_NOT U396 ( .A(n400), .Z(n399) );
  GTECH_NOT U397 ( .A(n389), .Z(n396) );
  GTECH_NAND2 U398 ( .A(I_b[1]), .B(I_a[2]), .Z(n389) );
  GTECH_NOT U399 ( .A(n387), .Z(n395) );
  GTECH_NAND2 U400 ( .A(I_b[0]), .B(I_a[3]), .Z(n387) );
  GTECH_NOT U401 ( .A(n376), .Z(n391) );
  GTECH_NAND3 U402 ( .A(I_a[0]), .B(n401), .C(I_b[2]), .Z(n376) );
  GTECH_XOR2 U403 ( .A(n402), .B(n401), .Z(N142) );
  GTECH_NOT U404 ( .A(n403), .Z(n401) );
  GTECH_XOR3 U405 ( .A(n397), .B(n398), .C(n400), .Z(n403) );
  GTECH_NAND3 U406 ( .A(n404), .B(I_b[0]), .C(I_a[1]), .Z(n400) );
  GTECH_NOT U407 ( .A(n405), .Z(n398) );
  GTECH_NAND2 U408 ( .A(I_a[1]), .B(I_b[1]), .Z(n405) );
  GTECH_NOT U409 ( .A(n406), .Z(n397) );
  GTECH_NAND2 U410 ( .A(I_b[0]), .B(I_a[2]), .Z(n406) );
  GTECH_AND2 U411 ( .A(I_b[2]), .B(I_a[0]), .Z(n402) );
  GTECH_XOR2 U412 ( .A(n404), .B(n407), .Z(N141) );
  GTECH_AND2 U413 ( .A(I_a[1]), .B(I_b[0]), .Z(n407) );
  GTECH_NOT U414 ( .A(n408), .Z(n404) );
  GTECH_NAND2 U415 ( .A(I_a[0]), .B(I_b[1]), .Z(n408) );
  GTECH_AND2 U416 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

