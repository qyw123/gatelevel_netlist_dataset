
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376;

  GTECH_MUX2 U135 ( .A(n274), .B(n275), .S(n276), .Z(sum[9]) );
  GTECH_OA21 U136 ( .A(n277), .B(n278), .C(n279), .Z(n276) );
  GTECH_OR_NOT U137 ( .A(n280), .B(n281), .Z(n275) );
  GTECH_XOR2 U138 ( .A(b[9]), .B(a[9]), .Z(n274) );
  GTECH_NAND2 U139 ( .A(n282), .B(n283), .Z(sum[8]) );
  GTECH_OAI21 U140 ( .A(n284), .B(n277), .C(n278), .Z(n282) );
  GTECH_MUX2 U141 ( .A(n285), .B(n286), .S(n287), .Z(sum[7]) );
  GTECH_XNOR2 U142 ( .A(n288), .B(n289), .Z(n286) );
  GTECH_XOR2 U143 ( .A(n288), .B(n290), .Z(n285) );
  GTECH_AND2 U144 ( .A(n291), .B(n292), .Z(n290) );
  GTECH_OAI21 U145 ( .A(b[6]), .B(a[6]), .C(n293), .Z(n292) );
  GTECH_XNOR2 U146 ( .A(a[7]), .B(b[7]), .Z(n288) );
  GTECH_OAI21 U147 ( .A(n294), .B(n291), .C(n295), .Z(sum[6]) );
  GTECH_MUX2 U148 ( .A(n296), .B(n297), .S(b[6]), .Z(n295) );
  GTECH_OR_NOT U149 ( .A(a[6]), .B(n294), .Z(n297) );
  GTECH_XOR2 U150 ( .A(a[6]), .B(n294), .Z(n296) );
  GTECH_AOI21 U151 ( .A(n287), .B(n298), .C(n293), .Z(n294) );
  GTECH_AOI21 U152 ( .A(n299), .B(n300), .C(n301), .Z(n293) );
  GTECH_MUX2 U153 ( .A(n302), .B(n303), .S(n304), .Z(sum[5]) );
  GTECH_AND2 U154 ( .A(n305), .B(n300), .Z(n304) );
  GTECH_OAI21 U155 ( .A(n306), .B(n287), .C(n307), .Z(n303) );
  GTECH_OAI21 U156 ( .A(n308), .B(n309), .C(n299), .Z(n302) );
  GTECH_NOT U157 ( .A(n307), .Z(n308) );
  GTECH_XOR2 U158 ( .A(n310), .B(n287), .Z(sum[4]) );
  GTECH_MUX2 U159 ( .A(n311), .B(n312), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U160 ( .A(n313), .B(n314), .Z(n312) );
  GTECH_XOR2 U161 ( .A(n315), .B(n313), .Z(n311) );
  GTECH_XOR2 U162 ( .A(a[3]), .B(b[3]), .Z(n313) );
  GTECH_ADD_ABC U163 ( .A(a[2]), .B(n316), .C(b[2]), .COUT(n315) );
  GTECH_MUX2 U164 ( .A(n317), .B(n318), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U165 ( .A(n319), .B(n320), .Z(n318) );
  GTECH_XOR2 U166 ( .A(n316), .B(n320), .Z(n317) );
  GTECH_XOR2 U167 ( .A(a[2]), .B(b[2]), .Z(n320) );
  GTECH_OA21 U168 ( .A(n321), .B(n322), .C(n323), .Z(n316) );
  GTECH_MUX2 U169 ( .A(n324), .B(n325), .S(n326), .Z(sum[1]) );
  GTECH_AND_NOT U170 ( .A(n323), .B(n321), .Z(n326) );
  GTECH_OAI21 U171 ( .A(cin), .B(n322), .C(n327), .Z(n325) );
  GTECH_AO21 U172 ( .A(n327), .B(cin), .C(n322), .Z(n324) );
  GTECH_MUX2 U173 ( .A(n328), .B(n329), .S(n330), .Z(sum[15]) );
  GTECH_XOR2 U174 ( .A(n331), .B(n332), .Z(n329) );
  GTECH_AOI21 U175 ( .A(n333), .B(n334), .C(n335), .Z(n332) );
  GTECH_XNOR2 U176 ( .A(n331), .B(n336), .Z(n328) );
  GTECH_XNOR2 U177 ( .A(a[15]), .B(b[15]), .Z(n331) );
  GTECH_MUX2 U178 ( .A(n337), .B(n338), .S(n339), .Z(sum[14]) );
  GTECH_AOI21 U179 ( .A(n340), .B(n341), .C(n334), .Z(n339) );
  GTECH_OA21 U180 ( .A(n342), .B(n343), .C(n344), .Z(n334) );
  GTECH_XOR2 U181 ( .A(b[14]), .B(a[14]), .Z(n338) );
  GTECH_OR_NOT U182 ( .A(n335), .B(n333), .Z(n337) );
  GTECH_MUX2 U183 ( .A(n345), .B(n346), .S(n347), .Z(sum[13]) );
  GTECH_OA21 U184 ( .A(n343), .B(n340), .C(n348), .Z(n347) );
  GTECH_OR_NOT U185 ( .A(n342), .B(n344), .Z(n346) );
  GTECH_XOR2 U186 ( .A(b[13]), .B(a[13]), .Z(n345) );
  GTECH_NAND2 U187 ( .A(n349), .B(n350), .Z(sum[12]) );
  GTECH_OAI21 U188 ( .A(n351), .B(n343), .C(n340), .Z(n349) );
  GTECH_MUX2 U189 ( .A(n352), .B(n353), .S(n354), .Z(sum[11]) );
  GTECH_XOR2 U190 ( .A(n355), .B(n356), .Z(n353) );
  GTECH_OA21 U191 ( .A(n357), .B(n358), .C(n359), .Z(n356) );
  GTECH_XNOR2 U192 ( .A(n355), .B(n360), .Z(n352) );
  GTECH_XNOR2 U193 ( .A(a[11]), .B(b[11]), .Z(n355) );
  GTECH_MUX2 U194 ( .A(n361), .B(n362), .S(n363), .Z(sum[10]) );
  GTECH_OA21 U195 ( .A(n354), .B(n364), .C(n358), .Z(n363) );
  GTECH_OAI21 U196 ( .A(n280), .B(n277), .C(n281), .Z(n358) );
  GTECH_XOR2 U197 ( .A(b[10]), .B(a[10]), .Z(n362) );
  GTECH_OR_NOT U198 ( .A(n357), .B(n359), .Z(n361) );
  GTECH_XNOR2 U199 ( .A(cin), .B(n365), .Z(sum[0]) );
  GTECH_OAI21 U200 ( .A(n330), .B(n366), .C(n350), .Z(cout) );
  GTECH_OR3 U201 ( .A(n351), .B(n343), .C(n340), .Z(n350) );
  GTECH_AND2 U202 ( .A(a[12]), .B(b[12]), .Z(n343) );
  GTECH_AOI21 U203 ( .A(n336), .B(a[15]), .C(n367), .Z(n366) );
  GTECH_OA21 U204 ( .A(a[15]), .B(n336), .C(b[15]), .Z(n367) );
  GTECH_AO21 U205 ( .A(n333), .B(n341), .C(n335), .Z(n336) );
  GTECH_AND2 U206 ( .A(a[14]), .B(b[14]), .Z(n335) );
  GTECH_OA21 U207 ( .A(n342), .B(n348), .C(n344), .Z(n341) );
  GTECH_OR2 U208 ( .A(b[13]), .B(a[13]), .Z(n344) );
  GTECH_NOT U209 ( .A(n351), .Z(n348) );
  GTECH_NOR2 U210 ( .A(b[12]), .B(a[12]), .Z(n351) );
  GTECH_AND2 U211 ( .A(a[13]), .B(b[13]), .Z(n342) );
  GTECH_OR2 U212 ( .A(a[14]), .B(b[14]), .Z(n333) );
  GTECH_NOT U213 ( .A(n340), .Z(n330) );
  GTECH_OAI21 U214 ( .A(n368), .B(n354), .C(n283), .Z(n340) );
  GTECH_OR3 U215 ( .A(n284), .B(n277), .C(n278), .Z(n283) );
  GTECH_AND2 U216 ( .A(b[8]), .B(a[8]), .Z(n277) );
  GTECH_NOT U217 ( .A(n278), .Z(n354) );
  GTECH_MUX2 U218 ( .A(n310), .B(n369), .S(n287), .Z(n278) );
  GTECH_NOT U219 ( .A(n309), .Z(n287) );
  GTECH_MUX2 U220 ( .A(n365), .B(n370), .S(cin), .Z(n309) );
  GTECH_AOI21 U221 ( .A(n314), .B(a[3]), .C(n371), .Z(n370) );
  GTECH_OA21 U222 ( .A(a[3]), .B(n314), .C(b[3]), .Z(n371) );
  GTECH_ADD_ABC U223 ( .A(n319), .B(a[2]), .C(b[2]), .COUT(n314) );
  GTECH_OA21 U224 ( .A(n321), .B(n327), .C(n323), .Z(n319) );
  GTECH_OR2 U225 ( .A(a[1]), .B(b[1]), .Z(n323) );
  GTECH_AND2 U226 ( .A(b[1]), .B(a[1]), .Z(n321) );
  GTECH_OR_NOT U227 ( .A(n322), .B(n327), .Z(n365) );
  GTECH_OR2 U228 ( .A(a[0]), .B(b[0]), .Z(n327) );
  GTECH_AND2 U229 ( .A(b[0]), .B(a[0]), .Z(n322) );
  GTECH_OA21 U230 ( .A(a[7]), .B(n289), .C(n372), .Z(n369) );
  GTECH_AO21 U231 ( .A(n289), .B(a[7]), .C(b[7]), .Z(n372) );
  GTECH_NAND2 U232 ( .A(n373), .B(n291), .Z(n289) );
  GTECH_NAND2 U233 ( .A(a[6]), .B(b[6]), .Z(n291) );
  GTECH_OAI21 U234 ( .A(a[6]), .B(b[6]), .C(n298), .Z(n373) );
  GTECH_OA21 U235 ( .A(n374), .B(n307), .C(n305), .Z(n298) );
  GTECH_NOT U236 ( .A(n301), .Z(n305) );
  GTECH_NOR2 U237 ( .A(b[5]), .B(a[5]), .Z(n301) );
  GTECH_NOT U238 ( .A(n300), .Z(n374) );
  GTECH_NAND2 U239 ( .A(a[5]), .B(b[5]), .Z(n300) );
  GTECH_AND_NOT U240 ( .A(n307), .B(n306), .Z(n310) );
  GTECH_NOT U241 ( .A(n299), .Z(n306) );
  GTECH_NAND2 U242 ( .A(b[4]), .B(a[4]), .Z(n299) );
  GTECH_OR2 U243 ( .A(a[4]), .B(b[4]), .Z(n307) );
  GTECH_AOI21 U244 ( .A(n360), .B(a[11]), .C(n375), .Z(n368) );
  GTECH_OA21 U245 ( .A(a[11]), .B(n360), .C(b[11]), .Z(n375) );
  GTECH_OAI21 U246 ( .A(n357), .B(n364), .C(n359), .Z(n360) );
  GTECH_NAND2 U247 ( .A(a[10]), .B(b[10]), .Z(n359) );
  GTECH_OAI21 U248 ( .A(n280), .B(n279), .C(n281), .Z(n364) );
  GTECH_OR_NOT U249 ( .A(a[9]), .B(n376), .Z(n281) );
  GTECH_NOT U250 ( .A(b[9]), .Z(n376) );
  GTECH_NOT U251 ( .A(n284), .Z(n279) );
  GTECH_NOR2 U252 ( .A(b[8]), .B(a[8]), .Z(n284) );
  GTECH_AND2 U253 ( .A(a[9]), .B(b[9]), .Z(n280) );
  GTECH_NOR2 U254 ( .A(b[10]), .B(a[10]), .Z(n357) );
endmodule

