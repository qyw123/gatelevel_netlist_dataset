
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390;

  GTECH_MUX2 U143 ( .A(n282), .B(n283), .S(n284), .Z(sum[9]) );
  GTECH_XNOR2 U144 ( .A(n285), .B(n286), .Z(n283) );
  GTECH_XNOR2 U145 ( .A(n285), .B(n287), .Z(n282) );
  GTECH_AOI21 U146 ( .A(a[9]), .B(b[9]), .C(n288), .Z(n285) );
  GTECH_NAND2 U147 ( .A(n289), .B(n290), .Z(sum[8]) );
  GTECH_OAI21 U148 ( .A(n291), .B(n286), .C(n284), .Z(n289) );
  GTECH_MUX2 U149 ( .A(n292), .B(n293), .S(n294), .Z(sum[7]) );
  GTECH_XOR2 U150 ( .A(n295), .B(n296), .Z(n293) );
  GTECH_XNOR2 U151 ( .A(n295), .B(n297), .Z(n292) );
  GTECH_AOI21 U152 ( .A(n298), .B(n299), .C(n300), .Z(n297) );
  GTECH_XOR2 U153 ( .A(a[7]), .B(b[7]), .Z(n295) );
  GTECH_MUX2 U154 ( .A(n301), .B(n302), .S(n303), .Z(sum[6]) );
  GTECH_AOI21 U155 ( .A(n294), .B(n304), .C(n299), .Z(n303) );
  GTECH_AOI21 U156 ( .A(n305), .B(n306), .C(n307), .Z(n299) );
  GTECH_XOR2 U157 ( .A(b[6]), .B(a[6]), .Z(n302) );
  GTECH_OR_NOT U158 ( .A(n300), .B(n298), .Z(n301) );
  GTECH_XOR2 U159 ( .A(n308), .B(n309), .Z(sum[5]) );
  GTECH_AOI21 U160 ( .A(n305), .B(n310), .C(n311), .Z(n309) );
  GTECH_AND_NOT U161 ( .A(n306), .B(n307), .Z(n308) );
  GTECH_XNOR2 U162 ( .A(n312), .B(n294), .Z(sum[4]) );
  GTECH_MUX2 U163 ( .A(n313), .B(n314), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U164 ( .A(n315), .B(n316), .Z(n314) );
  GTECH_XNOR2 U165 ( .A(n315), .B(n317), .Z(n313) );
  GTECH_AND2 U166 ( .A(n318), .B(n319), .Z(n317) );
  GTECH_OAI21 U167 ( .A(b[2]), .B(a[2]), .C(n320), .Z(n318) );
  GTECH_XOR2 U168 ( .A(a[3]), .B(b[3]), .Z(n315) );
  GTECH_MUX2 U169 ( .A(n321), .B(n322), .S(n323), .Z(sum[2]) );
  GTECH_NOT U170 ( .A(cin), .Z(n323) );
  GTECH_MUX2 U171 ( .A(n324), .B(n325), .S(n320), .Z(n322) );
  GTECH_OA21 U172 ( .A(n326), .B(n327), .C(n328), .Z(n320) );
  GTECH_MUX2 U173 ( .A(n324), .B(n325), .S(n329), .Z(n321) );
  GTECH_OAI21 U174 ( .A(b[2]), .B(a[2]), .C(n319), .Z(n325) );
  GTECH_XOR2 U175 ( .A(a[2]), .B(b[2]), .Z(n324) );
  GTECH_MUX2 U176 ( .A(n330), .B(n331), .S(n332), .Z(sum[1]) );
  GTECH_AND_NOT U177 ( .A(n328), .B(n327), .Z(n332) );
  GTECH_OAI21 U178 ( .A(cin), .B(n326), .C(n333), .Z(n331) );
  GTECH_AO21 U179 ( .A(n333), .B(cin), .C(n326), .Z(n330) );
  GTECH_AND_NOT U180 ( .A(a[0]), .B(n334), .Z(n326) );
  GTECH_MUX2 U181 ( .A(n335), .B(n336), .S(n337), .Z(sum[15]) );
  GTECH_XOR2 U182 ( .A(n338), .B(n339), .Z(n336) );
  GTECH_AND_NOT U183 ( .A(n340), .B(n341), .Z(n339) );
  GTECH_OAI21 U184 ( .A(b[14]), .B(a[14]), .C(n342), .Z(n340) );
  GTECH_XNOR2 U185 ( .A(n338), .B(n343), .Z(n335) );
  GTECH_XNOR2 U186 ( .A(a[15]), .B(b[15]), .Z(n338) );
  GTECH_AO21 U187 ( .A(n344), .B(n341), .C(n345), .Z(sum[14]) );
  GTECH_NOT U188 ( .A(n346), .Z(n345) );
  GTECH_MUX2 U189 ( .A(n347), .B(n348), .S(b[14]), .Z(n346) );
  GTECH_OR_NOT U190 ( .A(n344), .B(n349), .Z(n348) );
  GTECH_XOR2 U191 ( .A(n349), .B(n344), .Z(n347) );
  GTECH_NOT U192 ( .A(a[14]), .Z(n349) );
  GTECH_AO21 U193 ( .A(n350), .B(n351), .C(n342), .Z(n344) );
  GTECH_OA21 U194 ( .A(n352), .B(n353), .C(n354), .Z(n342) );
  GTECH_MUX2 U195 ( .A(n355), .B(n356), .S(n357), .Z(sum[13]) );
  GTECH_OA21 U196 ( .A(n353), .B(n350), .C(n358), .Z(n357) );
  GTECH_OR_NOT U197 ( .A(n352), .B(n354), .Z(n356) );
  GTECH_XNOR2 U198 ( .A(b[13]), .B(n359), .Z(n355) );
  GTECH_NAND2 U199 ( .A(n360), .B(n361), .Z(sum[12]) );
  GTECH_OAI21 U200 ( .A(n353), .B(n362), .C(n350), .Z(n360) );
  GTECH_MUX2 U201 ( .A(n363), .B(n364), .S(n284), .Z(sum[11]) );
  GTECH_XOR2 U202 ( .A(n365), .B(n366), .Z(n364) );
  GTECH_XNOR2 U203 ( .A(n365), .B(n367), .Z(n363) );
  GTECH_AND2 U204 ( .A(n368), .B(n369), .Z(n367) );
  GTECH_OAI21 U205 ( .A(b[10]), .B(a[10]), .C(n370), .Z(n368) );
  GTECH_XOR2 U206 ( .A(a[11]), .B(b[11]), .Z(n365) );
  GTECH_OAI21 U207 ( .A(n371), .B(n369), .C(n372), .Z(sum[10]) );
  GTECH_MUX2 U208 ( .A(n373), .B(n374), .S(b[10]), .Z(n372) );
  GTECH_OR_NOT U209 ( .A(a[10]), .B(n371), .Z(n374) );
  GTECH_XOR2 U210 ( .A(a[10]), .B(n371), .Z(n373) );
  GTECH_AOI21 U211 ( .A(n375), .B(n284), .C(n370), .Z(n371) );
  GTECH_OAI2N2 U212 ( .A(n288), .B(n287), .C(a[9]), .D(b[9]), .Z(n370) );
  GTECH_XNOR2 U213 ( .A(cin), .B(n376), .Z(sum[0]) );
  GTECH_OAI21 U214 ( .A(n337), .B(n377), .C(n361), .Z(cout) );
  GTECH_OR3 U215 ( .A(n353), .B(n362), .C(n350), .Z(n361) );
  GTECH_AND2 U216 ( .A(b[12]), .B(a[12]), .Z(n353) );
  GTECH_AOI21 U217 ( .A(n343), .B(a[15]), .C(n378), .Z(n377) );
  GTECH_OA21 U218 ( .A(a[15]), .B(n343), .C(b[15]), .Z(n378) );
  GTECH_OR_NOT U219 ( .A(n341), .B(n379), .Z(n343) );
  GTECH_OAI21 U220 ( .A(a[14]), .B(b[14]), .C(n351), .Z(n379) );
  GTECH_OA21 U221 ( .A(n352), .B(n358), .C(n354), .Z(n351) );
  GTECH_OR_NOT U222 ( .A(b[13]), .B(n359), .Z(n354) );
  GTECH_NOT U223 ( .A(a[13]), .Z(n359) );
  GTECH_NOT U224 ( .A(n362), .Z(n358) );
  GTECH_NOR2 U225 ( .A(b[12]), .B(a[12]), .Z(n362) );
  GTECH_AND2 U226 ( .A(b[13]), .B(a[13]), .Z(n352) );
  GTECH_AND2 U227 ( .A(b[14]), .B(a[14]), .Z(n341) );
  GTECH_NOT U228 ( .A(n350), .Z(n337) );
  GTECH_OAI21 U229 ( .A(n380), .B(n381), .C(n290), .Z(n350) );
  GTECH_OR3 U230 ( .A(n291), .B(n286), .C(n284), .Z(n290) );
  GTECH_NOT U231 ( .A(n381), .Z(n284) );
  GTECH_NOT U232 ( .A(n287), .Z(n291) );
  GTECH_NAND2 U233 ( .A(b[8]), .B(a[8]), .Z(n287) );
  GTECH_MUX2 U234 ( .A(n312), .B(n382), .S(n294), .Z(n381) );
  GTECH_NOT U235 ( .A(n310), .Z(n294) );
  GTECH_MUX2 U236 ( .A(n376), .B(n383), .S(cin), .Z(n310) );
  GTECH_AOI21 U237 ( .A(n316), .B(a[3]), .C(n384), .Z(n383) );
  GTECH_OA21 U238 ( .A(a[3]), .B(n316), .C(b[3]), .Z(n384) );
  GTECH_NAND2 U239 ( .A(n319), .B(n385), .Z(n316) );
  GTECH_OAI21 U240 ( .A(a[2]), .B(b[2]), .C(n329), .Z(n385) );
  GTECH_OA21 U241 ( .A(n327), .B(n333), .C(n328), .Z(n329) );
  GTECH_OR_NOT U242 ( .A(a[1]), .B(n386), .Z(n328) );
  GTECH_OR_NOT U243 ( .A(a[0]), .B(n334), .Z(n333) );
  GTECH_NOT U244 ( .A(b[0]), .Z(n334) );
  GTECH_AND_NOT U245 ( .A(a[1]), .B(n386), .Z(n327) );
  GTECH_NOT U246 ( .A(b[1]), .Z(n386) );
  GTECH_NAND2 U247 ( .A(b[2]), .B(a[2]), .Z(n319) );
  GTECH_XNOR2 U248 ( .A(a[0]), .B(b[0]), .Z(n376) );
  GTECH_AOI21 U249 ( .A(n296), .B(a[7]), .C(n387), .Z(n382) );
  GTECH_OA21 U250 ( .A(a[7]), .B(n296), .C(b[7]), .Z(n387) );
  GTECH_AO21 U251 ( .A(n298), .B(n304), .C(n300), .Z(n296) );
  GTECH_AND_NOT U252 ( .A(b[6]), .B(n388), .Z(n300) );
  GTECH_AOI21 U253 ( .A(n306), .B(n311), .C(n307), .Z(n304) );
  GTECH_NOR2 U254 ( .A(a[5]), .B(b[5]), .Z(n307) );
  GTECH_NAND2 U255 ( .A(a[5]), .B(b[5]), .Z(n306) );
  GTECH_OR_NOT U256 ( .A(b[6]), .B(n388), .Z(n298) );
  GTECH_NOT U257 ( .A(a[6]), .Z(n388) );
  GTECH_OR_NOT U258 ( .A(n311), .B(n305), .Z(n312) );
  GTECH_NAND2 U259 ( .A(a[4]), .B(b[4]), .Z(n305) );
  GTECH_NOR2 U260 ( .A(b[4]), .B(a[4]), .Z(n311) );
  GTECH_AOI21 U261 ( .A(n366), .B(a[11]), .C(n389), .Z(n380) );
  GTECH_OA21 U262 ( .A(a[11]), .B(n366), .C(b[11]), .Z(n389) );
  GTECH_NAND2 U263 ( .A(n390), .B(n369), .Z(n366) );
  GTECH_NAND2 U264 ( .A(a[10]), .B(b[10]), .Z(n369) );
  GTECH_OAI21 U265 ( .A(a[10]), .B(b[10]), .C(n375), .Z(n390) );
  GTECH_OAI2N2 U266 ( .A(n286), .B(n288), .C(a[9]), .D(b[9]), .Z(n375) );
  GTECH_NOR2 U267 ( .A(a[9]), .B(b[9]), .Z(n288) );
  GTECH_NOR2 U268 ( .A(b[8]), .B(a[8]), .Z(n286) );
endmodule

