
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NAND2 U83 ( .A(n93), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI21 U86 ( .A(n98), .B(n99), .C(n100), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_NAND2 U88 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U89 ( .A(n104), .Z(n84) );
  GTECH_NAND2 U90 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_XOR2 U91 ( .A(n106), .B(n105), .Z(N153) );
  GTECH_NOT U92 ( .A(n107), .Z(n105) );
  GTECH_XNOR3 U93 ( .A(n108), .B(n93), .C(n109), .Z(n107) );
  GTECH_NOT U94 ( .A(n95), .Z(n109) );
  GTECH_XNOR3 U95 ( .A(n101), .B(n103), .C(n98), .Z(n95) );
  GTECH_NOT U96 ( .A(n102), .Z(n98) );
  GTECH_OAI21 U97 ( .A(n110), .B(n111), .C(n112), .Z(n102) );
  GTECH_OAI21 U98 ( .A(n113), .B(n114), .C(n115), .Z(n112) );
  GTECH_NOT U99 ( .A(n116), .Z(n103) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n116) );
  GTECH_NOT U101 ( .A(n99), .Z(n101) );
  GTECH_NAND2 U102 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U103 ( .A(n117), .B(n118), .C(n119), .COUT(n93) );
  GTECH_NOT U104 ( .A(n120), .Z(n119) );
  GTECH_XOR2 U105 ( .A(n121), .B(n122), .Z(n118) );
  GTECH_AND2 U106 ( .A(I_a[7]), .B(I_b[5]), .Z(n122) );
  GTECH_NOT U107 ( .A(n94), .Z(n108) );
  GTECH_NAND2 U108 ( .A(I_a[7]), .B(n123), .Z(n94) );
  GTECH_NOT U109 ( .A(n124), .Z(n106) );
  GTECH_NAND2 U110 ( .A(n125), .B(n126), .Z(n124) );
  GTECH_NOT U111 ( .A(n127), .Z(n126) );
  GTECH_XOR2 U112 ( .A(n127), .B(n128), .Z(N152) );
  GTECH_NOT U113 ( .A(n125), .Z(n128) );
  GTECH_XOR4 U114 ( .A(n129), .B(n121), .C(n120), .D(n117), .Z(n125) );
  GTECH_ADD_ABC U115 ( .A(n130), .B(n131), .C(n132), .COUT(n117) );
  GTECH_XNOR3 U116 ( .A(n133), .B(n134), .C(n135), .Z(n131) );
  GTECH_XNOR3 U117 ( .A(n113), .B(n115), .C(n110), .Z(n120) );
  GTECH_NOT U118 ( .A(n114), .Z(n110) );
  GTECH_OAI21 U119 ( .A(n136), .B(n137), .C(n138), .Z(n114) );
  GTECH_OAI21 U120 ( .A(n139), .B(n140), .C(n141), .Z(n138) );
  GTECH_NOT U121 ( .A(n142), .Z(n115) );
  GTECH_NAND2 U122 ( .A(I_b[7]), .B(I_a[5]), .Z(n142) );
  GTECH_NOT U123 ( .A(n111), .Z(n113) );
  GTECH_NAND2 U124 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_NOT U125 ( .A(n123), .Z(n121) );
  GTECH_OAI21 U126 ( .A(n143), .B(n144), .C(n145), .Z(n123) );
  GTECH_OAI21 U127 ( .A(n133), .B(n135), .C(n134), .Z(n145) );
  GTECH_AND2 U128 ( .A(I_a[7]), .B(I_b[5]), .Z(n129) );
  GTECH_ADD_ABC U129 ( .A(n146), .B(n147), .C(n148), .COUT(n127) );
  GTECH_OA22 U130 ( .A(n149), .B(n150), .C(n151), .D(n152), .Z(n147) );
  GTECH_OA21 U131 ( .A(n153), .B(n154), .C(n155), .Z(n146) );
  GTECH_XNOR3 U132 ( .A(n156), .B(n148), .C(n157), .Z(N151) );
  GTECH_OA21 U133 ( .A(n153), .B(n154), .C(n155), .Z(n157) );
  GTECH_OAI21 U134 ( .A(n158), .B(n159), .C(n160), .Z(n155) );
  GTECH_XOR2 U135 ( .A(n130), .B(n161), .Z(n148) );
  GTECH_XOR4 U136 ( .A(n134), .B(n143), .C(n132), .D(n133), .Z(n161) );
  GTECH_NOT U137 ( .A(n144), .Z(n133) );
  GTECH_NAND2 U138 ( .A(I_a[7]), .B(I_b[4]), .Z(n144) );
  GTECH_NOT U139 ( .A(n162), .Z(n132) );
  GTECH_XNOR3 U140 ( .A(n139), .B(n141), .C(n136), .Z(n162) );
  GTECH_NOT U141 ( .A(n140), .Z(n136) );
  GTECH_OAI21 U142 ( .A(n163), .B(n164), .C(n165), .Z(n140) );
  GTECH_OAI21 U143 ( .A(n166), .B(n167), .C(n168), .Z(n165) );
  GTECH_NOT U144 ( .A(n169), .Z(n141) );
  GTECH_NAND2 U145 ( .A(I_b[7]), .B(I_a[4]), .Z(n169) );
  GTECH_NOT U146 ( .A(n137), .Z(n139) );
  GTECH_NAND2 U147 ( .A(I_b[6]), .B(I_a[5]), .Z(n137) );
  GTECH_NOT U148 ( .A(n135), .Z(n143) );
  GTECH_OAI21 U149 ( .A(n170), .B(n171), .C(n172), .Z(n135) );
  GTECH_OAI21 U150 ( .A(n173), .B(n174), .C(n175), .Z(n172) );
  GTECH_NOT U151 ( .A(n176), .Z(n134) );
  GTECH_NAND2 U152 ( .A(I_a[6]), .B(I_b[5]), .Z(n176) );
  GTECH_ADD_ABC U153 ( .A(n177), .B(n178), .C(n179), .COUT(n130) );
  GTECH_NOT U154 ( .A(n180), .Z(n179) );
  GTECH_XNOR3 U155 ( .A(n173), .B(n175), .C(n174), .Z(n178) );
  GTECH_OA22 U156 ( .A(n149), .B(n150), .C(n151), .D(n152), .Z(n156) );
  GTECH_NOT U157 ( .A(n181), .Z(n152) );
  GTECH_NOT U158 ( .A(I_a[7]), .Z(n150) );
  GTECH_XNOR3 U159 ( .A(n153), .B(n158), .C(n160), .Z(N150) );
  GTECH_XOR2 U160 ( .A(n182), .B(n177), .Z(n160) );
  GTECH_ADD_ABC U161 ( .A(n183), .B(n184), .C(n185), .COUT(n177) );
  GTECH_NOT U162 ( .A(n186), .Z(n185) );
  GTECH_XNOR3 U163 ( .A(n187), .B(n188), .C(n189), .Z(n184) );
  GTECH_XOR4 U164 ( .A(n175), .B(n170), .C(n180), .D(n173), .Z(n182) );
  GTECH_NOT U165 ( .A(n171), .Z(n173) );
  GTECH_NAND2 U166 ( .A(I_a[6]), .B(I_b[4]), .Z(n171) );
  GTECH_XNOR3 U167 ( .A(n166), .B(n168), .C(n163), .Z(n180) );
  GTECH_NOT U168 ( .A(n167), .Z(n163) );
  GTECH_OAI21 U169 ( .A(n190), .B(n191), .C(n192), .Z(n167) );
  GTECH_OAI21 U170 ( .A(n193), .B(n194), .C(n195), .Z(n192) );
  GTECH_NOT U171 ( .A(n196), .Z(n168) );
  GTECH_NAND2 U172 ( .A(I_b[7]), .B(I_a[3]), .Z(n196) );
  GTECH_NOT U173 ( .A(n164), .Z(n166) );
  GTECH_NAND2 U174 ( .A(I_b[6]), .B(I_a[4]), .Z(n164) );
  GTECH_NOT U175 ( .A(n174), .Z(n170) );
  GTECH_OAI21 U176 ( .A(n197), .B(n198), .C(n199), .Z(n174) );
  GTECH_OAI21 U177 ( .A(n187), .B(n189), .C(n188), .Z(n199) );
  GTECH_NOT U178 ( .A(n200), .Z(n175) );
  GTECH_NAND2 U179 ( .A(I_a[5]), .B(I_b[5]), .Z(n200) );
  GTECH_NOT U180 ( .A(n154), .Z(n158) );
  GTECH_XOR2 U181 ( .A(n181), .B(n151), .Z(n154) );
  GTECH_NOT U182 ( .A(n201), .Z(n151) );
  GTECH_OAI2N2 U183 ( .A(n202), .B(n203), .C(n204), .D(n205), .Z(n201) );
  GTECH_NAND2 U184 ( .A(n202), .B(n203), .Z(n205) );
  GTECH_XOR2 U185 ( .A(n206), .B(n149), .Z(n181) );
  GTECH_OA21 U186 ( .A(n207), .B(n208), .C(n209), .Z(n149) );
  GTECH_OAI21 U187 ( .A(n210), .B(n211), .C(n212), .Z(n209) );
  GTECH_NAND2 U188 ( .A(I_a[7]), .B(I_b[3]), .Z(n206) );
  GTECH_NOT U189 ( .A(n159), .Z(n153) );
  GTECH_OAI2N2 U190 ( .A(n213), .B(n214), .C(n215), .D(n216), .Z(n159) );
  GTECH_NAND2 U191 ( .A(n213), .B(n214), .Z(n216) );
  GTECH_XNOR3 U192 ( .A(n213), .B(n217), .C(n215), .Z(N149) );
  GTECH_XOR2 U193 ( .A(n218), .B(n183), .Z(n215) );
  GTECH_ADD_ABC U194 ( .A(n219), .B(n220), .C(n221), .COUT(n183) );
  GTECH_XNOR3 U195 ( .A(n222), .B(n223), .C(n224), .Z(n220) );
  GTECH_OA21 U196 ( .A(n225), .B(n226), .C(n227), .Z(n219) );
  GTECH_XOR4 U197 ( .A(n188), .B(n197), .C(n186), .D(n187), .Z(n218) );
  GTECH_NOT U198 ( .A(n198), .Z(n187) );
  GTECH_NAND2 U199 ( .A(I_a[5]), .B(I_b[4]), .Z(n198) );
  GTECH_XNOR3 U200 ( .A(n193), .B(n195), .C(n190), .Z(n186) );
  GTECH_NOT U201 ( .A(n194), .Z(n190) );
  GTECH_OAI21 U202 ( .A(n228), .B(n229), .C(n230), .Z(n194) );
  GTECH_NOT U203 ( .A(n231), .Z(n195) );
  GTECH_NAND2 U204 ( .A(I_b[7]), .B(I_a[2]), .Z(n231) );
  GTECH_NOT U205 ( .A(n191), .Z(n193) );
  GTECH_NAND2 U206 ( .A(I_b[6]), .B(I_a[3]), .Z(n191) );
  GTECH_NOT U207 ( .A(n189), .Z(n197) );
  GTECH_OAI21 U208 ( .A(n232), .B(n233), .C(n234), .Z(n189) );
  GTECH_OAI21 U209 ( .A(n222), .B(n224), .C(n223), .Z(n234) );
  GTECH_NOT U210 ( .A(n235), .Z(n188) );
  GTECH_NAND2 U211 ( .A(I_b[5]), .B(I_a[4]), .Z(n235) );
  GTECH_NOT U212 ( .A(n214), .Z(n217) );
  GTECH_XNOR3 U213 ( .A(n236), .B(n202), .C(n237), .Z(n214) );
  GTECH_NOT U214 ( .A(n204), .Z(n237) );
  GTECH_XNOR3 U215 ( .A(n210), .B(n212), .C(n207), .Z(n204) );
  GTECH_NOT U216 ( .A(n211), .Z(n207) );
  GTECH_OAI21 U217 ( .A(n238), .B(n239), .C(n240), .Z(n211) );
  GTECH_OAI21 U218 ( .A(n241), .B(n242), .C(n243), .Z(n240) );
  GTECH_NOT U219 ( .A(n244), .Z(n212) );
  GTECH_NAND2 U220 ( .A(I_a[6]), .B(I_b[3]), .Z(n244) );
  GTECH_NOT U221 ( .A(n208), .Z(n210) );
  GTECH_NAND2 U222 ( .A(I_a[7]), .B(I_b[2]), .Z(n208) );
  GTECH_ADD_ABC U223 ( .A(n245), .B(n246), .C(n247), .COUT(n202) );
  GTECH_NOT U224 ( .A(n248), .Z(n247) );
  GTECH_XOR2 U225 ( .A(n249), .B(n250), .Z(n246) );
  GTECH_AND2 U226 ( .A(I_a[7]), .B(I_b[1]), .Z(n250) );
  GTECH_NOT U227 ( .A(n203), .Z(n236) );
  GTECH_NAND2 U228 ( .A(I_a[7]), .B(n251), .Z(n203) );
  GTECH_ADD_ABC U229 ( .A(n252), .B(n253), .C(n254), .COUT(n213) );
  GTECH_XNOR3 U230 ( .A(n245), .B(n255), .C(n248), .Z(n253) );
  GTECH_XOR2 U231 ( .A(n256), .B(n252), .Z(N148) );
  GTECH_ADD_ABC U232 ( .A(n257), .B(n258), .C(n259), .COUT(n252) );
  GTECH_NOT U233 ( .A(n260), .Z(n259) );
  GTECH_XNOR3 U234 ( .A(n261), .B(n262), .C(n263), .Z(n258) );
  GTECH_XOR4 U235 ( .A(n255), .B(n245), .C(n248), .D(n254), .Z(n256) );
  GTECH_XOR2 U236 ( .A(n264), .B(n265), .Z(n254) );
  GTECH_XOR4 U237 ( .A(n223), .B(n232), .C(n221), .D(n222), .Z(n265) );
  GTECH_NOT U238 ( .A(n233), .Z(n222) );
  GTECH_NAND2 U239 ( .A(I_b[4]), .B(I_a[4]), .Z(n233) );
  GTECH_XNOR3 U240 ( .A(n266), .B(n267), .C(n268), .Z(n221) );
  GTECH_NOT U241 ( .A(n230), .Z(n268) );
  GTECH_NAND3 U242 ( .A(I_b[6]), .B(I_a[1]), .C(n269), .Z(n230) );
  GTECH_NOT U243 ( .A(n229), .Z(n267) );
  GTECH_NAND2 U244 ( .A(I_b[7]), .B(I_a[1]), .Z(n229) );
  GTECH_NOT U245 ( .A(n228), .Z(n266) );
  GTECH_NAND2 U246 ( .A(I_b[6]), .B(I_a[2]), .Z(n228) );
  GTECH_NOT U247 ( .A(n224), .Z(n232) );
  GTECH_OAI21 U248 ( .A(n270), .B(n271), .C(n272), .Z(n224) );
  GTECH_OAI21 U249 ( .A(n273), .B(n274), .C(n275), .Z(n272) );
  GTECH_NOT U250 ( .A(n276), .Z(n223) );
  GTECH_NAND2 U251 ( .A(I_b[5]), .B(I_a[3]), .Z(n276) );
  GTECH_OA21 U252 ( .A(n225), .B(n226), .C(n227), .Z(n264) );
  GTECH_OAI21 U253 ( .A(n277), .B(n278), .C(n279), .Z(n227) );
  GTECH_XNOR3 U254 ( .A(n241), .B(n243), .C(n238), .Z(n248) );
  GTECH_NOT U255 ( .A(n242), .Z(n238) );
  GTECH_OAI21 U256 ( .A(n280), .B(n281), .C(n282), .Z(n242) );
  GTECH_OAI21 U257 ( .A(n283), .B(n284), .C(n285), .Z(n282) );
  GTECH_NOT U258 ( .A(n286), .Z(n243) );
  GTECH_NAND2 U259 ( .A(I_a[5]), .B(I_b[3]), .Z(n286) );
  GTECH_NOT U260 ( .A(n239), .Z(n241) );
  GTECH_NAND2 U261 ( .A(I_a[6]), .B(I_b[2]), .Z(n239) );
  GTECH_ADD_ABC U262 ( .A(n261), .B(n287), .C(n288), .COUT(n245) );
  GTECH_XNOR3 U263 ( .A(n289), .B(n290), .C(n291), .Z(n287) );
  GTECH_XOR2 U264 ( .A(n292), .B(n249), .Z(n255) );
  GTECH_NOT U265 ( .A(n251), .Z(n249) );
  GTECH_OAI21 U266 ( .A(n293), .B(n294), .C(n295), .Z(n251) );
  GTECH_OAI21 U267 ( .A(n289), .B(n291), .C(n290), .Z(n295) );
  GTECH_AND2 U268 ( .A(I_a[7]), .B(I_b[1]), .Z(n292) );
  GTECH_XOR2 U269 ( .A(n296), .B(n257), .Z(N147) );
  GTECH_ADD_ABC U270 ( .A(n297), .B(n298), .C(n299), .COUT(n257) );
  GTECH_XNOR3 U271 ( .A(n300), .B(n301), .C(n302), .Z(n298) );
  GTECH_OA21 U272 ( .A(n303), .B(n304), .C(n305), .Z(n297) );
  GTECH_XOR4 U273 ( .A(n262), .B(n288), .C(n260), .D(n261), .Z(n296) );
  GTECH_ADD_ABC U274 ( .A(n300), .B(n306), .C(n307), .COUT(n261) );
  GTECH_NOT U275 ( .A(n302), .Z(n307) );
  GTECH_XNOR3 U276 ( .A(n308), .B(n309), .C(n310), .Z(n306) );
  GTECH_XNOR3 U277 ( .A(n279), .B(n226), .C(n278), .Z(n260) );
  GTECH_NOT U278 ( .A(n225), .Z(n278) );
  GTECH_XOR2 U279 ( .A(n311), .B(n269), .Z(n225) );
  GTECH_NOT U280 ( .A(n312), .Z(n269) );
  GTECH_NAND2 U281 ( .A(I_b[7]), .B(I_a[0]), .Z(n312) );
  GTECH_NAND2 U282 ( .A(I_b[6]), .B(I_a[1]), .Z(n311) );
  GTECH_NOT U283 ( .A(n277), .Z(n226) );
  GTECH_XNOR3 U284 ( .A(n273), .B(n275), .C(n270), .Z(n277) );
  GTECH_NOT U285 ( .A(n274), .Z(n270) );
  GTECH_OAI21 U286 ( .A(n313), .B(n314), .C(n315), .Z(n274) );
  GTECH_NOT U287 ( .A(n316), .Z(n275) );
  GTECH_NAND2 U288 ( .A(I_b[5]), .B(I_a[2]), .Z(n316) );
  GTECH_NOT U289 ( .A(n271), .Z(n273) );
  GTECH_NAND2 U290 ( .A(I_b[4]), .B(I_a[3]), .Z(n271) );
  GTECH_NOT U291 ( .A(n317), .Z(n279) );
  GTECH_NAND3 U292 ( .A(I_a[0]), .B(n318), .C(I_b[6]), .Z(n317) );
  GTECH_NOT U293 ( .A(n319), .Z(n318) );
  GTECH_NOT U294 ( .A(n263), .Z(n288) );
  GTECH_XNOR3 U295 ( .A(n283), .B(n285), .C(n280), .Z(n263) );
  GTECH_NOT U296 ( .A(n284), .Z(n280) );
  GTECH_OAI21 U297 ( .A(n320), .B(n321), .C(n322), .Z(n284) );
  GTECH_OAI21 U298 ( .A(n323), .B(n324), .C(n325), .Z(n322) );
  GTECH_NOT U299 ( .A(n326), .Z(n285) );
  GTECH_NAND2 U300 ( .A(I_b[3]), .B(I_a[4]), .Z(n326) );
  GTECH_NOT U301 ( .A(n281), .Z(n283) );
  GTECH_NAND2 U302 ( .A(I_a[5]), .B(I_b[2]), .Z(n281) );
  GTECH_NOT U303 ( .A(n327), .Z(n262) );
  GTECH_XNOR3 U304 ( .A(n289), .B(n290), .C(n293), .Z(n327) );
  GTECH_NOT U305 ( .A(n291), .Z(n293) );
  GTECH_OAI21 U306 ( .A(n328), .B(n329), .C(n330), .Z(n291) );
  GTECH_OAI21 U307 ( .A(n308), .B(n310), .C(n309), .Z(n330) );
  GTECH_NOT U308 ( .A(n331), .Z(n290) );
  GTECH_NAND2 U309 ( .A(I_a[6]), .B(I_b[1]), .Z(n331) );
  GTECH_NOT U310 ( .A(n294), .Z(n289) );
  GTECH_NAND2 U311 ( .A(I_a[7]), .B(I_b[0]), .Z(n294) );
  GTECH_XOR2 U312 ( .A(n332), .B(n333), .Z(N146) );
  GTECH_OA21 U313 ( .A(n303), .B(n304), .C(n305), .Z(n333) );
  GTECH_OAI21 U314 ( .A(n334), .B(n335), .C(n336), .Z(n305) );
  GTECH_XOR4 U315 ( .A(n301), .B(n300), .C(n302), .D(n299), .Z(n332) );
  GTECH_XOR2 U316 ( .A(n319), .B(n337), .Z(n299) );
  GTECH_AND2 U317 ( .A(I_b[6]), .B(I_a[0]), .Z(n337) );
  GTECH_XNOR3 U318 ( .A(n338), .B(n339), .C(n340), .Z(n319) );
  GTECH_NOT U319 ( .A(n315), .Z(n340) );
  GTECH_NAND3 U320 ( .A(I_b[4]), .B(I_a[1]), .C(n341), .Z(n315) );
  GTECH_NOT U321 ( .A(n314), .Z(n339) );
  GTECH_NAND2 U322 ( .A(I_b[5]), .B(I_a[1]), .Z(n314) );
  GTECH_NOT U323 ( .A(n313), .Z(n338) );
  GTECH_NAND2 U324 ( .A(I_b[4]), .B(I_a[2]), .Z(n313) );
  GTECH_XNOR3 U325 ( .A(n323), .B(n325), .C(n320), .Z(n302) );
  GTECH_NOT U326 ( .A(n324), .Z(n320) );
  GTECH_OAI21 U327 ( .A(n342), .B(n343), .C(n344), .Z(n324) );
  GTECH_OAI21 U328 ( .A(n345), .B(n346), .C(n347), .Z(n344) );
  GTECH_NOT U329 ( .A(n348), .Z(n325) );
  GTECH_NAND2 U330 ( .A(I_b[3]), .B(I_a[3]), .Z(n348) );
  GTECH_NOT U331 ( .A(n321), .Z(n323) );
  GTECH_NAND2 U332 ( .A(I_b[2]), .B(I_a[4]), .Z(n321) );
  GTECH_ADD_ABC U333 ( .A(n349), .B(n350), .C(n351), .COUT(n300) );
  GTECH_NOT U334 ( .A(n352), .Z(n351) );
  GTECH_XNOR3 U335 ( .A(n353), .B(n354), .C(n355), .Z(n350) );
  GTECH_NOT U336 ( .A(n356), .Z(n301) );
  GTECH_XNOR3 U337 ( .A(n308), .B(n309), .C(n328), .Z(n356) );
  GTECH_NOT U338 ( .A(n310), .Z(n328) );
  GTECH_OAI21 U339 ( .A(n357), .B(n358), .C(n359), .Z(n310) );
  GTECH_OAI21 U340 ( .A(n353), .B(n355), .C(n354), .Z(n359) );
  GTECH_NOT U341 ( .A(n360), .Z(n309) );
  GTECH_NAND2 U342 ( .A(I_a[5]), .B(I_b[1]), .Z(n360) );
  GTECH_NOT U343 ( .A(n329), .Z(n308) );
  GTECH_NAND2 U344 ( .A(I_a[6]), .B(I_b[0]), .Z(n329) );
  GTECH_XNOR3 U345 ( .A(n336), .B(n304), .C(n335), .Z(N145) );
  GTECH_NOT U346 ( .A(n303), .Z(n335) );
  GTECH_XOR2 U347 ( .A(n361), .B(n341), .Z(n303) );
  GTECH_NOT U348 ( .A(n362), .Z(n341) );
  GTECH_NAND2 U349 ( .A(I_b[5]), .B(I_a[0]), .Z(n362) );
  GTECH_NAND2 U350 ( .A(I_b[4]), .B(I_a[1]), .Z(n361) );
  GTECH_NOT U351 ( .A(n334), .Z(n304) );
  GTECH_XOR2 U352 ( .A(n363), .B(n349), .Z(n334) );
  GTECH_ADD_ABC U353 ( .A(n364), .B(n365), .C(n366), .COUT(n349) );
  GTECH_XNOR3 U354 ( .A(n367), .B(n368), .C(n369), .Z(n365) );
  GTECH_OA21 U355 ( .A(n370), .B(n371), .C(n372), .Z(n364) );
  GTECH_XOR4 U356 ( .A(n354), .B(n357), .C(n352), .D(n353), .Z(n363) );
  GTECH_NOT U357 ( .A(n358), .Z(n353) );
  GTECH_NAND2 U358 ( .A(I_a[5]), .B(I_b[0]), .Z(n358) );
  GTECH_XNOR3 U359 ( .A(n345), .B(n347), .C(n342), .Z(n352) );
  GTECH_NOT U360 ( .A(n346), .Z(n342) );
  GTECH_OAI21 U361 ( .A(n373), .B(n374), .C(n375), .Z(n346) );
  GTECH_NOT U362 ( .A(n376), .Z(n347) );
  GTECH_NAND2 U363 ( .A(I_b[3]), .B(I_a[2]), .Z(n376) );
  GTECH_NOT U364 ( .A(n343), .Z(n345) );
  GTECH_NAND2 U365 ( .A(I_b[2]), .B(I_a[3]), .Z(n343) );
  GTECH_NOT U366 ( .A(n355), .Z(n357) );
  GTECH_OAI21 U367 ( .A(n377), .B(n378), .C(n379), .Z(n355) );
  GTECH_OAI21 U368 ( .A(n367), .B(n369), .C(n368), .Z(n379) );
  GTECH_NOT U369 ( .A(n378), .Z(n367) );
  GTECH_NOT U370 ( .A(n380), .Z(n354) );
  GTECH_NAND2 U371 ( .A(I_a[4]), .B(I_b[1]), .Z(n380) );
  GTECH_NOT U372 ( .A(n381), .Z(n336) );
  GTECH_NAND3 U373 ( .A(I_a[0]), .B(n382), .C(I_b[4]), .Z(n381) );
  GTECH_XOR2 U374 ( .A(n383), .B(n382), .Z(N144) );
  GTECH_XOR2 U375 ( .A(n384), .B(n385), .Z(n382) );
  GTECH_OA21 U376 ( .A(n370), .B(n371), .C(n372), .Z(n385) );
  GTECH_OAI21 U377 ( .A(n386), .B(n387), .C(n388), .Z(n372) );
  GTECH_XOR4 U378 ( .A(n368), .B(n377), .C(n378), .D(n366), .Z(n384) );
  GTECH_XNOR3 U379 ( .A(n389), .B(n390), .C(n391), .Z(n366) );
  GTECH_NOT U380 ( .A(n375), .Z(n391) );
  GTECH_NAND3 U381 ( .A(I_b[2]), .B(I_a[1]), .C(n392), .Z(n375) );
  GTECH_NOT U382 ( .A(n374), .Z(n390) );
  GTECH_NAND2 U383 ( .A(I_b[3]), .B(I_a[1]), .Z(n374) );
  GTECH_NOT U384 ( .A(n373), .Z(n389) );
  GTECH_NAND2 U385 ( .A(I_b[2]), .B(I_a[2]), .Z(n373) );
  GTECH_NAND2 U386 ( .A(I_a[4]), .B(I_b[0]), .Z(n378) );
  GTECH_NOT U387 ( .A(n369), .Z(n377) );
  GTECH_OAI21 U388 ( .A(n393), .B(n394), .C(n395), .Z(n369) );
  GTECH_OAI21 U389 ( .A(n396), .B(n397), .C(n398), .Z(n395) );
  GTECH_NOT U390 ( .A(n399), .Z(n368) );
  GTECH_NAND2 U391 ( .A(I_a[3]), .B(I_b[1]), .Z(n399) );
  GTECH_AND2 U392 ( .A(I_b[4]), .B(I_a[0]), .Z(n383) );
  GTECH_XNOR3 U393 ( .A(n388), .B(n371), .C(n387), .Z(N143) );
  GTECH_NOT U394 ( .A(n370), .Z(n387) );
  GTECH_XOR2 U395 ( .A(n400), .B(n392), .Z(n370) );
  GTECH_NOT U396 ( .A(n401), .Z(n392) );
  GTECH_NAND2 U397 ( .A(I_b[3]), .B(I_a[0]), .Z(n401) );
  GTECH_NAND2 U398 ( .A(I_b[2]), .B(I_a[1]), .Z(n400) );
  GTECH_NOT U399 ( .A(n386), .Z(n371) );
  GTECH_XNOR3 U400 ( .A(n396), .B(n398), .C(n393), .Z(n386) );
  GTECH_NOT U401 ( .A(n397), .Z(n393) );
  GTECH_OAI21 U402 ( .A(n402), .B(n403), .C(n404), .Z(n397) );
  GTECH_NOT U403 ( .A(n405), .Z(n398) );
  GTECH_NAND2 U404 ( .A(I_b[1]), .B(I_a[2]), .Z(n405) );
  GTECH_NOT U405 ( .A(n394), .Z(n396) );
  GTECH_NAND2 U406 ( .A(I_b[0]), .B(I_a[3]), .Z(n394) );
  GTECH_NOT U407 ( .A(n406), .Z(n388) );
  GTECH_NAND3 U408 ( .A(I_a[0]), .B(n407), .C(I_b[2]), .Z(n406) );
  GTECH_XOR2 U409 ( .A(n408), .B(n407), .Z(N142) );
  GTECH_NOT U410 ( .A(n409), .Z(n407) );
  GTECH_XNOR3 U411 ( .A(n410), .B(n411), .C(n412), .Z(n409) );
  GTECH_NOT U412 ( .A(n404), .Z(n412) );
  GTECH_NAND3 U413 ( .A(n413), .B(I_b[0]), .C(I_a[1]), .Z(n404) );
  GTECH_NOT U414 ( .A(n402), .Z(n411) );
  GTECH_NAND2 U415 ( .A(I_a[1]), .B(I_b[1]), .Z(n402) );
  GTECH_NOT U416 ( .A(n403), .Z(n410) );
  GTECH_NAND2 U417 ( .A(I_b[0]), .B(I_a[2]), .Z(n403) );
  GTECH_AND2 U418 ( .A(I_b[2]), .B(I_a[0]), .Z(n408) );
  GTECH_XOR2 U419 ( .A(n413), .B(n414), .Z(N141) );
  GTECH_AND2 U420 ( .A(I_a[1]), .B(I_b[0]), .Z(n414) );
  GTECH_NOT U421 ( .A(n415), .Z(n413) );
  GTECH_NAND2 U422 ( .A(I_a[0]), .B(I_b[1]), .Z(n415) );
  GTECH_AND2 U423 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

