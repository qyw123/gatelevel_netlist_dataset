
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374;

  GTECH_MUX2 U127 ( .A(n266), .B(n267), .S(n268), .Z(sum[9]) );
  GTECH_XNOR2 U128 ( .A(n269), .B(n270), .Z(n267) );
  GTECH_XNOR2 U129 ( .A(n271), .B(n269), .Z(n266) );
  GTECH_OR_NOT U130 ( .A(n272), .B(n273), .Z(n269) );
  GTECH_XNOR2 U131 ( .A(n274), .B(n275), .Z(sum[8]) );
  GTECH_MUX2 U132 ( .A(n276), .B(n277), .S(n278), .Z(sum[7]) );
  GTECH_XNOR2 U133 ( .A(n279), .B(n280), .Z(n277) );
  GTECH_AOI21 U134 ( .A(n281), .B(n282), .C(n283), .Z(n280) );
  GTECH_XNOR2 U135 ( .A(n279), .B(n284), .Z(n276) );
  GTECH_XOR2 U136 ( .A(a[7]), .B(b[7]), .Z(n279) );
  GTECH_MUX2 U137 ( .A(n285), .B(n286), .S(n278), .Z(sum[6]) );
  GTECH_XOR2 U138 ( .A(n287), .B(n282), .Z(n286) );
  GTECH_OR_NOT U139 ( .A(n288), .B(n289), .Z(n282) );
  GTECH_OR3 U140 ( .A(n290), .B(n291), .C(n292), .Z(n289) );
  GTECH_XOR2 U141 ( .A(n287), .B(n293), .Z(n285) );
  GTECH_AND_NOT U142 ( .A(n281), .B(n283), .Z(n287) );
  GTECH_XOR2 U143 ( .A(n294), .B(n295), .Z(sum[5]) );
  GTECH_OA22 U144 ( .A(n278), .B(n292), .C(n296), .D(n290), .Z(n295) );
  GTECH_AND_NOT U145 ( .A(n292), .B(n297), .Z(n296) );
  GTECH_NOT U146 ( .A(n278), .Z(n297) );
  GTECH_OR2 U147 ( .A(n288), .B(n291), .Z(n294) );
  GTECH_XOR2 U148 ( .A(n298), .B(n278), .Z(sum[4]) );
  GTECH_MUX2 U149 ( .A(n299), .B(n300), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U150 ( .A(n301), .B(n302), .Z(n300) );
  GTECH_XNOR2 U151 ( .A(n301), .B(n303), .Z(n299) );
  GTECH_OA21 U152 ( .A(n304), .B(n305), .C(n306), .Z(n303) );
  GTECH_XOR2 U153 ( .A(a[3]), .B(b[3]), .Z(n301) );
  GTECH_MUX2 U154 ( .A(n307), .B(n308), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U155 ( .A(n309), .B(n310), .Z(n308) );
  GTECH_XNOR2 U156 ( .A(n309), .B(n305), .Z(n307) );
  GTECH_AOI21 U157 ( .A(n311), .B(n312), .C(n313), .Z(n305) );
  GTECH_AND_NOT U158 ( .A(n306), .B(n304), .Z(n309) );
  GTECH_NOT U159 ( .A(n314), .Z(sum[1]) );
  GTECH_MUX2 U160 ( .A(n315), .B(n316), .S(n317), .Z(n314) );
  GTECH_AND_NOT U161 ( .A(n311), .B(n313), .Z(n317) );
  GTECH_OA21 U162 ( .A(cin), .B(n312), .C(n318), .Z(n316) );
  GTECH_AOI21 U163 ( .A(n318), .B(cin), .C(n312), .Z(n315) );
  GTECH_MUX2 U164 ( .A(n319), .B(n320), .S(n321), .Z(sum[15]) );
  GTECH_XNOR2 U165 ( .A(n322), .B(n323), .Z(n320) );
  GTECH_AOI21 U166 ( .A(n324), .B(n325), .C(n326), .Z(n323) );
  GTECH_XNOR2 U167 ( .A(n322), .B(n327), .Z(n319) );
  GTECH_XNOR2 U168 ( .A(n328), .B(b[15]), .Z(n322) );
  GTECH_MUX2 U169 ( .A(n329), .B(n330), .S(n321), .Z(sum[14]) );
  GTECH_XNOR2 U170 ( .A(n325), .B(n331), .Z(n330) );
  GTECH_OA21 U171 ( .A(n332), .B(n333), .C(n334), .Z(n325) );
  GTECH_XNOR2 U172 ( .A(n335), .B(n331), .Z(n329) );
  GTECH_OR_NOT U173 ( .A(n326), .B(n324), .Z(n331) );
  GTECH_MUX2 U174 ( .A(n336), .B(n337), .S(n321), .Z(sum[13]) );
  GTECH_XOR2 U175 ( .A(n333), .B(n338), .Z(n337) );
  GTECH_XOR2 U176 ( .A(n338), .B(n339), .Z(n336) );
  GTECH_AOI21 U177 ( .A(n340), .B(n341), .C(n332), .Z(n338) );
  GTECH_OR_NOT U178 ( .A(n342), .B(n343), .Z(sum[12]) );
  GTECH_OA21 U179 ( .A(n333), .B(n344), .C(n345), .Z(n342) );
  GTECH_MUX2 U180 ( .A(n346), .B(n347), .S(n268), .Z(sum[11]) );
  GTECH_XOR2 U181 ( .A(n348), .B(n349), .Z(n347) );
  GTECH_XOR2 U182 ( .A(n348), .B(n350), .Z(n346) );
  GTECH_OA21 U183 ( .A(n351), .B(n352), .C(n353), .Z(n350) );
  GTECH_XOR2 U184 ( .A(n354), .B(b[11]), .Z(n348) );
  GTECH_MUX2 U185 ( .A(n355), .B(n356), .S(n275), .Z(sum[10]) );
  GTECH_XNOR2 U186 ( .A(n357), .B(n352), .Z(n356) );
  GTECH_AOI21 U187 ( .A(n273), .B(n271), .C(n272), .Z(n352) );
  GTECH_XNOR2 U188 ( .A(n357), .B(n358), .Z(n355) );
  GTECH_AND_NOT U189 ( .A(n353), .B(n351), .Z(n357) );
  GTECH_OR_NOT U190 ( .A(n359), .B(n360), .Z(sum[0]) );
  GTECH_OA21 U191 ( .A(n361), .B(n312), .C(cin), .Z(n359) );
  GTECH_NOT U192 ( .A(n362), .Z(cout) );
  GTECH_OA21 U193 ( .A(n363), .B(n321), .C(n343), .Z(n362) );
  GTECH_OR3 U194 ( .A(n333), .B(n344), .C(n345), .Z(n343) );
  GTECH_AND2 U195 ( .A(a[12]), .B(b[12]), .Z(n333) );
  GTECH_NOT U196 ( .A(n345), .Z(n321) );
  GTECH_MUX2 U197 ( .A(n274), .B(n364), .S(n268), .Z(n345) );
  GTECH_NOT U198 ( .A(n275), .Z(n268) );
  GTECH_MUX2 U199 ( .A(n365), .B(n298), .S(n278), .Z(n275) );
  GTECH_OA21 U200 ( .A(n366), .B(n367), .C(n360), .Z(n278) );
  GTECH_OR3 U201 ( .A(n312), .B(cin), .C(n361), .Z(n360) );
  GTECH_AND2 U202 ( .A(b[0]), .B(a[0]), .Z(n312) );
  GTECH_NOT U203 ( .A(cin), .Z(n367) );
  GTECH_AOI2N2 U204 ( .A(n368), .B(b[3]), .C(n302), .D(n369), .Z(n366) );
  GTECH_NAND2 U205 ( .A(n369), .B(n302), .Z(n368) );
  GTECH_OA21 U206 ( .A(n304), .B(n310), .C(n306), .Z(n302) );
  GTECH_NAND2 U207 ( .A(a[2]), .B(b[2]), .Z(n306) );
  GTECH_AOI21 U208 ( .A(n311), .B(n318), .C(n313), .Z(n310) );
  GTECH_AND2 U209 ( .A(a[1]), .B(b[1]), .Z(n313) );
  GTECH_NOT U210 ( .A(n361), .Z(n318) );
  GTECH_NOR2 U211 ( .A(a[0]), .B(b[0]), .Z(n361) );
  GTECH_OR2 U212 ( .A(a[1]), .B(b[1]), .Z(n311) );
  GTECH_NOR2 U213 ( .A(b[2]), .B(a[2]), .Z(n304) );
  GTECH_NOT U214 ( .A(a[3]), .Z(n369) );
  GTECH_XNOR2 U215 ( .A(a[4]), .B(b[4]), .Z(n298) );
  GTECH_AOI2N2 U216 ( .A(n370), .B(b[7]), .C(n284), .D(n371), .Z(n365) );
  GTECH_NAND2 U217 ( .A(n371), .B(n284), .Z(n370) );
  GTECH_AOI21 U218 ( .A(n281), .B(n293), .C(n283), .Z(n284) );
  GTECH_AND2 U219 ( .A(b[6]), .B(a[6]), .Z(n283) );
  GTECH_OR2 U220 ( .A(n372), .B(n288), .Z(n293) );
  GTECH_AND2 U221 ( .A(b[5]), .B(a[5]), .Z(n288) );
  GTECH_AOI21 U222 ( .A(n290), .B(n292), .C(n291), .Z(n372) );
  GTECH_NOR2 U223 ( .A(b[5]), .B(a[5]), .Z(n291) );
  GTECH_NOT U224 ( .A(a[4]), .Z(n292) );
  GTECH_NOT U225 ( .A(b[4]), .Z(n290) );
  GTECH_OR2 U226 ( .A(b[6]), .B(a[6]), .Z(n281) );
  GTECH_NOT U227 ( .A(a[7]), .Z(n371) );
  GTECH_AOI2N2 U228 ( .A(n354), .B(n349), .C(b[11]), .D(n373), .Z(n364) );
  GTECH_NOR2 U229 ( .A(n354), .B(n349), .Z(n373) );
  GTECH_OA21 U230 ( .A(n351), .B(n358), .C(n353), .Z(n349) );
  GTECH_NAND2 U231 ( .A(a[10]), .B(b[10]), .Z(n353) );
  GTECH_AOI21 U232 ( .A(n273), .B(n270), .C(n272), .Z(n358) );
  GTECH_AND2 U233 ( .A(b[9]), .B(a[9]), .Z(n272) );
  GTECH_OR2 U234 ( .A(b[9]), .B(a[9]), .Z(n273) );
  GTECH_NOR2 U235 ( .A(b[10]), .B(a[10]), .Z(n351) );
  GTECH_NOT U236 ( .A(a[11]), .Z(n354) );
  GTECH_AND_NOT U237 ( .A(n270), .B(n271), .Z(n274) );
  GTECH_AND2 U238 ( .A(b[8]), .B(a[8]), .Z(n271) );
  GTECH_OR2 U239 ( .A(a[8]), .B(b[8]), .Z(n270) );
  GTECH_AOI2N2 U240 ( .A(n374), .B(b[15]), .C(n327), .D(n328), .Z(n363) );
  GTECH_NAND2 U241 ( .A(n328), .B(n327), .Z(n374) );
  GTECH_AOI21 U242 ( .A(n324), .B(n335), .C(n326), .Z(n327) );
  GTECH_AND2 U243 ( .A(b[14]), .B(a[14]), .Z(n326) );
  GTECH_OA21 U244 ( .A(n332), .B(n339), .C(n334), .Z(n335) );
  GTECH_NAND2 U245 ( .A(n341), .B(n340), .Z(n334) );
  GTECH_NOT U246 ( .A(a[13]), .Z(n340) );
  GTECH_NOT U247 ( .A(b[13]), .Z(n341) );
  GTECH_NOT U248 ( .A(n344), .Z(n339) );
  GTECH_NOR2 U249 ( .A(b[12]), .B(a[12]), .Z(n344) );
  GTECH_AND2 U250 ( .A(a[13]), .B(b[13]), .Z(n332) );
  GTECH_OR2 U251 ( .A(b[14]), .B(a[14]), .Z(n324) );
  GTECH_NOT U252 ( .A(a[15]), .Z(n328) );
endmodule

