
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382;

  GTECH_MUX2 U130 ( .A(n269), .B(n270), .S(n271), .Z(sum[9]) );
  GTECH_XNOR2 U131 ( .A(n272), .B(n273), .Z(n270) );
  GTECH_XOR2 U132 ( .A(n274), .B(n273), .Z(n269) );
  GTECH_AO21 U133 ( .A(n275), .B(n276), .C(n277), .Z(n273) );
  GTECH_OR_NOT U134 ( .A(n278), .B(n279), .Z(sum[8]) );
  GTECH_AO21 U135 ( .A(n272), .B(n274), .C(n280), .Z(n279) );
  GTECH_MUX2 U136 ( .A(n281), .B(n282), .S(n283), .Z(sum[7]) );
  GTECH_XOR2 U137 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_XOR2 U138 ( .A(n286), .B(n284), .Z(n281) );
  GTECH_XOR2 U139 ( .A(a[7]), .B(b[7]), .Z(n284) );
  GTECH_OA22 U140 ( .A(a[6]), .B(n287), .C(b[6]), .D(n288), .Z(n286) );
  GTECH_AND2 U141 ( .A(n287), .B(a[6]), .Z(n288) );
  GTECH_MUX2 U142 ( .A(n289), .B(n290), .S(n283), .Z(sum[6]) );
  GTECH_XNOR2 U143 ( .A(n291), .B(n292), .Z(n290) );
  GTECH_XNOR2 U144 ( .A(n291), .B(n287), .Z(n289) );
  GTECH_AO21 U145 ( .A(n293), .B(n294), .C(n295), .Z(n287) );
  GTECH_XNOR2 U146 ( .A(a[6]), .B(b[6]), .Z(n291) );
  GTECH_MUX2 U147 ( .A(n296), .B(n297), .S(n298), .Z(sum[5]) );
  GTECH_AND_NOT U148 ( .A(n294), .B(n295), .Z(n298) );
  GTECH_AO21 U149 ( .A(n299), .B(n300), .C(n301), .Z(n297) );
  GTECH_OAI22 U150 ( .A(n302), .B(n303), .C(n299), .D(n304), .Z(n296) );
  GTECH_NOT U151 ( .A(n283), .Z(n299) );
  GTECH_AND_NOT U152 ( .A(n304), .B(n283), .Z(n302) );
  GTECH_XOR2 U153 ( .A(n283), .B(n305), .Z(sum[4]) );
  GTECH_MUX2 U154 ( .A(n306), .B(n307), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U155 ( .A(n308), .B(n309), .Z(n307) );
  GTECH_XNOR2 U156 ( .A(n310), .B(n308), .Z(n306) );
  GTECH_XNOR2 U157 ( .A(a[3]), .B(b[3]), .Z(n308) );
  GTECH_OA22 U158 ( .A(a[2]), .B(n311), .C(b[2]), .D(n312), .Z(n310) );
  GTECH_AND2 U159 ( .A(n311), .B(a[2]), .Z(n312) );
  GTECH_MUX2 U160 ( .A(n313), .B(n314), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U161 ( .A(n315), .B(n316), .Z(n314) );
  GTECH_XNOR2 U162 ( .A(n315), .B(n311), .Z(n313) );
  GTECH_AO21 U163 ( .A(n317), .B(n318), .C(n319), .Z(n311) );
  GTECH_XNOR2 U164 ( .A(a[2]), .B(b[2]), .Z(n315) );
  GTECH_MUX2 U165 ( .A(n320), .B(n321), .S(cin), .Z(sum[1]) );
  GTECH_XNOR2 U166 ( .A(n322), .B(n323), .Z(n321) );
  GTECH_XNOR2 U167 ( .A(n317), .B(n322), .Z(n320) );
  GTECH_OR_NOT U168 ( .A(n319), .B(n318), .Z(n322) );
  GTECH_MUX2 U169 ( .A(n324), .B(n325), .S(n326), .Z(sum[15]) );
  GTECH_XNOR2 U170 ( .A(n327), .B(n328), .Z(n325) );
  GTECH_XOR2 U171 ( .A(n329), .B(n327), .Z(n324) );
  GTECH_XOR2 U172 ( .A(a[15]), .B(b[15]), .Z(n327) );
  GTECH_OA22 U173 ( .A(a[14]), .B(n330), .C(b[14]), .D(n331), .Z(n329) );
  GTECH_AND_NOT U174 ( .A(n330), .B(n332), .Z(n331) );
  GTECH_MUX2 U175 ( .A(n333), .B(n334), .S(n326), .Z(sum[14]) );
  GTECH_XOR2 U176 ( .A(n335), .B(n336), .Z(n334) );
  GTECH_XNOR2 U177 ( .A(n335), .B(n330), .Z(n333) );
  GTECH_AO21 U178 ( .A(n337), .B(n338), .C(n339), .Z(n330) );
  GTECH_XNOR2 U179 ( .A(n332), .B(n340), .Z(n335) );
  GTECH_MUX2 U180 ( .A(n341), .B(n342), .S(n326), .Z(sum[13]) );
  GTECH_XNOR2 U181 ( .A(n343), .B(n344), .Z(n342) );
  GTECH_XNOR2 U182 ( .A(n337), .B(n343), .Z(n341) );
  GTECH_OR_NOT U183 ( .A(n339), .B(n338), .Z(n343) );
  GTECH_OR_NOT U184 ( .A(n345), .B(n346), .Z(sum[12]) );
  GTECH_AO21 U185 ( .A(n344), .B(n347), .C(n348), .Z(n346) );
  GTECH_MUX2 U186 ( .A(n349), .B(n350), .S(n271), .Z(sum[11]) );
  GTECH_XOR2 U187 ( .A(n351), .B(n352), .Z(n350) );
  GTECH_XOR2 U188 ( .A(n353), .B(n351), .Z(n349) );
  GTECH_XNOR2 U189 ( .A(a[11]), .B(n354), .Z(n351) );
  GTECH_ADD_ABC U190 ( .A(a[10]), .B(n355), .C(b[10]), .COUT(n353) );
  GTECH_MUX2 U191 ( .A(n356), .B(n357), .S(n271), .Z(sum[10]) );
  GTECH_XOR2 U192 ( .A(n358), .B(n359), .Z(n357) );
  GTECH_XOR2 U193 ( .A(n355), .B(n359), .Z(n356) );
  GTECH_XOR2 U194 ( .A(a[10]), .B(b[10]), .Z(n359) );
  GTECH_AOI21 U195 ( .A(n274), .B(n360), .C(n361), .Z(n355) );
  GTECH_XOR2 U196 ( .A(cin), .B(n362), .Z(sum[0]) );
  GTECH_AO21 U197 ( .A(n363), .B(n326), .C(n345), .Z(cout) );
  GTECH_AND3 U198 ( .A(n344), .B(n347), .C(n348), .Z(n345) );
  GTECH_NOT U199 ( .A(n337), .Z(n347) );
  GTECH_AND2 U200 ( .A(b[12]), .B(a[12]), .Z(n337) );
  GTECH_NOT U201 ( .A(n348), .Z(n326) );
  GTECH_AOI21 U202 ( .A(n271), .B(n364), .C(n278), .Z(n348) );
  GTECH_AND3 U203 ( .A(n272), .B(n274), .C(n280), .Z(n278) );
  GTECH_NOT U204 ( .A(n271), .Z(n280) );
  GTECH_NAND2 U205 ( .A(b[8]), .B(a[8]), .Z(n274) );
  GTECH_OAI22 U206 ( .A(n365), .B(n354), .C(n366), .D(n367), .Z(n364) );
  GTECH_NOT U207 ( .A(n352), .Z(n366) );
  GTECH_NOT U208 ( .A(b[11]), .Z(n354) );
  GTECH_AND_NOT U209 ( .A(n367), .B(n352), .Z(n365) );
  GTECH_ADD_ABC U210 ( .A(n358), .B(a[10]), .C(b[10]), .COUT(n352) );
  GTECH_AOI21 U211 ( .A(n368), .B(n360), .C(n361), .Z(n358) );
  GTECH_AND_NOT U212 ( .A(n275), .B(a[9]), .Z(n361) );
  GTECH_NOT U213 ( .A(n277), .Z(n360) );
  GTECH_NOR2 U214 ( .A(n276), .B(n275), .Z(n277) );
  GTECH_NOT U215 ( .A(b[9]), .Z(n275) );
  GTECH_NOT U216 ( .A(a[9]), .Z(n276) );
  GTECH_NOT U217 ( .A(n272), .Z(n368) );
  GTECH_OR2 U218 ( .A(a[8]), .B(b[8]), .Z(n272) );
  GTECH_NOT U219 ( .A(a[11]), .Z(n367) );
  GTECH_MUX2 U220 ( .A(n305), .B(n369), .S(n283), .Z(n271) );
  GTECH_MUX2 U221 ( .A(n362), .B(n370), .S(cin), .Z(n283) );
  GTECH_OA22 U222 ( .A(a[3]), .B(n309), .C(b[3]), .D(n371), .Z(n370) );
  GTECH_AND2 U223 ( .A(n309), .B(a[3]), .Z(n371) );
  GTECH_OAI2N2 U224 ( .A(n372), .B(n373), .C(n316), .D(a[2]), .Z(n309) );
  GTECH_NOT U225 ( .A(n374), .Z(n316) );
  GTECH_NOT U226 ( .A(b[2]), .Z(n373) );
  GTECH_AND_NOT U227 ( .A(n374), .B(a[2]), .Z(n372) );
  GTECH_AOI21 U228 ( .A(n318), .B(n323), .C(n319), .Z(n374) );
  GTECH_AND2 U229 ( .A(a[1]), .B(b[1]), .Z(n319) );
  GTECH_OR2 U230 ( .A(b[1]), .B(a[1]), .Z(n318) );
  GTECH_AND_NOT U231 ( .A(n323), .B(n317), .Z(n362) );
  GTECH_AND2 U232 ( .A(a[0]), .B(b[0]), .Z(n317) );
  GTECH_OR2 U233 ( .A(b[0]), .B(a[0]), .Z(n323) );
  GTECH_OA22 U234 ( .A(a[7]), .B(n285), .C(b[7]), .D(n375), .Z(n369) );
  GTECH_AND2 U235 ( .A(n285), .B(a[7]), .Z(n375) );
  GTECH_OAI2N2 U236 ( .A(n376), .B(n377), .C(n292), .D(a[6]), .Z(n285) );
  GTECH_NOT U237 ( .A(n378), .Z(n292) );
  GTECH_NOT U238 ( .A(b[6]), .Z(n377) );
  GTECH_AND_NOT U239 ( .A(n378), .B(a[6]), .Z(n376) );
  GTECH_AOI21 U240 ( .A(n379), .B(n294), .C(n295), .Z(n378) );
  GTECH_AND2 U241 ( .A(a[5]), .B(b[5]), .Z(n295) );
  GTECH_OR2 U242 ( .A(b[5]), .B(a[5]), .Z(n294) );
  GTECH_AND2 U243 ( .A(n379), .B(n300), .Z(n305) );
  GTECH_NOT U244 ( .A(n293), .Z(n300) );
  GTECH_NOR2 U245 ( .A(n303), .B(n304), .Z(n293) );
  GTECH_NOT U246 ( .A(a[4]), .Z(n304) );
  GTECH_NOT U247 ( .A(b[4]), .Z(n303) );
  GTECH_NOT U248 ( .A(n301), .Z(n379) );
  GTECH_NOR2 U249 ( .A(b[4]), .B(a[4]), .Z(n301) );
  GTECH_AO22 U250 ( .A(n380), .B(a[15]), .C(n381), .D(b[15]), .Z(n363) );
  GTECH_OR_NOT U251 ( .A(a[15]), .B(n328), .Z(n381) );
  GTECH_NOT U252 ( .A(n328), .Z(n380) );
  GTECH_OA22 U253 ( .A(n336), .B(n332), .C(n382), .D(n340), .Z(n328) );
  GTECH_NOT U254 ( .A(b[14]), .Z(n340) );
  GTECH_AND_NOT U255 ( .A(n336), .B(a[14]), .Z(n382) );
  GTECH_NOT U256 ( .A(a[14]), .Z(n332) );
  GTECH_AOI21 U257 ( .A(n344), .B(n338), .C(n339), .Z(n336) );
  GTECH_AND2 U258 ( .A(a[13]), .B(b[13]), .Z(n339) );
  GTECH_OR2 U259 ( .A(b[13]), .B(a[13]), .Z(n338) );
  GTECH_OR2 U260 ( .A(a[12]), .B(b[12]), .Z(n344) );
endmodule

