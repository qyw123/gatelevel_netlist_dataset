
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n115, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n115), .K(n115), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n252) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n115), .K(n115), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n115), .K(n115), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n115), .K(n115), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n115), .K(n115), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n115), .K(n115), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]) );
  GTECH_FJK1S A_reg_15_ ( .J(n115), .K(n115), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n268) );
  GTECH_FJK1S A_reg_14_ ( .J(n115), .K(n115), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n267) );
  GTECH_FJK1S A_reg_13_ ( .J(n115), .K(n115), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n266) );
  GTECH_FJK1S A_reg_12_ ( .J(n115), .K(n115), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n265) );
  GTECH_FJK1S A_reg_11_ ( .J(n115), .K(n115), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n264) );
  GTECH_FJK1S A_reg_10_ ( .J(n115), .K(n115), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n263) );
  GTECH_FJK1S A_reg_9_ ( .J(n115), .K(n115), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n262) );
  GTECH_FJK1S A_reg_8_ ( .J(n115), .K(n115), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n261) );
  GTECH_FJK1S A_reg_7_ ( .J(n115), .K(n115), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n260) );
  GTECH_FJK1S A_reg_6_ ( .J(n115), .K(n115), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n259) );
  GTECH_FJK1S A_reg_5_ ( .J(n115), .K(n115), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n258) );
  GTECH_FJK1S A_reg_4_ ( .J(n115), .K(n115), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n257) );
  GTECH_FJK1S A_reg_3_ ( .J(n115), .K(n115), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n256) );
  GTECH_FJK1S A_reg_2_ ( .J(n115), .K(n115), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n255) );
  GTECH_FJK1S A_reg_1_ ( .J(n115), .K(n115), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n254) );
  GTECH_FJK1S A_reg_0_ ( .J(n115), .K(n115), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n253) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n115), .K(n115), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n115), .K(n115), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n115), .K(n115), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n115), .K(n115), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n115), .K(n115), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n115), .K(n115), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n115), .K(n115), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n115), .K(n115), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n115), .K(n115), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n115), .K(n115), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n115), .K(n115), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n115), .K(n115), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n115), .K(n115), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n115), .K(n115), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n115), .K(n115), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n115), .K(n115), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n115), .K(n115), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n115), .K(n115), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n115), .K(n115), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n115), .K(n115), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n115), .K(n115), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n115), .K(n115), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n115), .K(n115), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n115), .K(n115), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n115), .K(n115), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n115), .K(n115), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n115), .K(n115), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n115), .K(n115), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n115), .K(n115), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n115), .K(n115), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n115), .K(n115), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n115), .K(n115), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n115), .K(n115), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n115), .K(n115), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n115), .K(n115), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n115), .K(n115), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n115), .K(n115), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n115), .K(n115), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n115), .K(n115), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n115), .K(n115), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n115), .K(n115), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n115), .K(n115), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n115), .K(n115), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n115), .K(n115), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n115), .K(n115), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n115), .K(n115), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n115), .K(n115), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n115), .K(n115), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n115), .K(n115), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n115), .K(n115), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n115), .K(n115), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n115), .K(n115), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n115), .K(n115), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n115), .K(n115), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n115), .K(n115), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n115), .K(n115), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n115), .K(n115), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n115), .K(n115), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n115), .K(n115), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n115), .K(n115), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n115), .K(n115), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n115), .K(n115), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n115), .K(n115), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n115), .K(n115), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n115), .K(n115), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n115), .K(n115), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U254 ( .Z(n115) );
  GTECH_NOT U255 ( .A(n270), .Z(N99) );
  GTECH_AOI222 U256 ( .A(n271), .B(n272), .C(n273), .D(n274), .E(n275), .F(
        n276), .Z(n270) );
  GTECH_NOT U257 ( .A(n277), .Z(N98) );
  GTECH_AOI222 U258 ( .A(n273), .B(n278), .C(n279), .D(n280), .E(R[15]), .F(
        n281), .Z(n277) );
  GTECH_OR_NOT U259 ( .A(n275), .B(n282), .Z(n279) );
  GTECH_OAI2N2 U260 ( .A(n13), .B(n283), .C(R[14]), .D(n281), .Z(N97) );
  GTECH_OAI2N2 U261 ( .A(n14), .B(n283), .C(R[13]), .D(n281), .Z(N96) );
  GTECH_OAI2N2 U262 ( .A(n15), .B(n283), .C(R[12]), .D(n281), .Z(N95) );
  GTECH_OAI2N2 U263 ( .A(n16), .B(n283), .C(R[11]), .D(n281), .Z(N94) );
  GTECH_OAI2N2 U264 ( .A(n17), .B(n283), .C(R[10]), .D(n281), .Z(N93) );
  GTECH_OAI2N2 U265 ( .A(n18), .B(n283), .C(R[9]), .D(n281), .Z(N92) );
  GTECH_OAI2N2 U266 ( .A(n19), .B(n283), .C(R[8]), .D(n281), .Z(N91) );
  GTECH_OAI2N2 U267 ( .A(n20), .B(n283), .C(R[7]), .D(n281), .Z(N90) );
  GTECH_OAI2N2 U268 ( .A(n21), .B(n283), .C(R[6]), .D(n281), .Z(N89) );
  GTECH_OAI2N2 U269 ( .A(n22), .B(n283), .C(R[5]), .D(n281), .Z(N88) );
  GTECH_OAI2N2 U270 ( .A(n23), .B(n283), .C(R[4]), .D(n281), .Z(N87) );
  GTECH_OAI2N2 U271 ( .A(n24), .B(n283), .C(R[3]), .D(n281), .Z(N86) );
  GTECH_OAI2N2 U272 ( .A(n25), .B(n283), .C(R[2]), .D(n281), .Z(N85) );
  GTECH_OAI2N2 U273 ( .A(n26), .B(n283), .C(R[1]), .D(n281), .Z(N84) );
  GTECH_OAI2N2 U274 ( .A(n27), .B(n283), .C(R[0]), .D(n281), .Z(N83) );
  GTECH_AND2 U275 ( .A(M[15]), .B(n281), .Z(N42) );
  GTECH_AND2 U276 ( .A(M[14]), .B(n281), .Z(N39) );
  GTECH_AND2 U277 ( .A(M[13]), .B(n281), .Z(N38) );
  GTECH_AND2 U278 ( .A(M[12]), .B(n281), .Z(N37) );
  GTECH_AND2 U279 ( .A(M[11]), .B(n281), .Z(N36) );
  GTECH_AND2 U280 ( .A(M[10]), .B(n281), .Z(N35) );
  GTECH_AND2 U281 ( .A(M[9]), .B(n281), .Z(N34) );
  GTECH_AND2 U282 ( .A(M[8]), .B(n281), .Z(N33) );
  GTECH_AND2 U283 ( .A(M[7]), .B(n281), .Z(N32) );
  GTECH_AND2 U284 ( .A(M[6]), .B(n281), .Z(N31) );
  GTECH_AND2 U285 ( .A(M[5]), .B(n281), .Z(N30) );
  GTECH_AND2 U286 ( .A(M[4]), .B(n281), .Z(N29) );
  GTECH_AND2 U287 ( .A(M[3]), .B(n281), .Z(N28) );
  GTECH_AND2 U288 ( .A(M[2]), .B(n281), .Z(N27) );
  GTECH_AND2 U289 ( .A(M[1]), .B(n281), .Z(N26) );
  GTECH_AND2 U290 ( .A(M[0]), .B(n281), .Z(N25) );
  GTECH_OAI21 U291 ( .A(n283), .B(n284), .C(n285), .Z(N19) );
  GTECH_OR_NOT U292 ( .A(n9), .B(n286), .Z(n284) );
  GTECH_OR3 U293 ( .A(Rst), .B(Ld), .C(n287), .Z(N18) );
  GTECH_AOI21 U294 ( .A(n286), .B(n288), .C(n283), .Z(N17) );
  GTECH_OR_NOT U295 ( .A(n8), .B(n289), .Z(n288) );
  GTECH_AOI21 U296 ( .A(n289), .B(n290), .C(n283), .Z(N16) );
  GTECH_OR_NOT U297 ( .A(n7), .B(n291), .Z(n290) );
  GTECH_NOT U298 ( .A(n292), .Z(N152) );
  GTECH_AOI222 U299 ( .A(n293), .B(n294), .C(n295), .D(n296), .E(n297), .F(
        n298), .Z(n292) );
  GTECH_OR_NOT U300 ( .A(N155), .B(n299), .Z(N151) );
  GTECH_NOT U301 ( .A(n300), .Z(N150) );
  GTECH_AOI222 U302 ( .A(n301), .B(n293), .C(n295), .D(n302), .E(n297), .F(
        n303), .Z(n300) );
  GTECH_MUX2 U303 ( .A(n304), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND2 U304 ( .A(n287), .B(n305), .Z(n304) );
  GTECH_NOT U305 ( .A(n306), .Z(N149) );
  GTECH_AOI222 U306 ( .A(n307), .B(n293), .C(n295), .D(n308), .E(n297), .F(
        n309), .Z(n306) );
  GTECH_NOT U307 ( .A(n310), .Z(N148) );
  GTECH_AOI222 U308 ( .A(n311), .B(n293), .C(n295), .D(n312), .E(n297), .F(
        n313), .Z(n310) );
  GTECH_NOT U309 ( .A(n314), .Z(N147) );
  GTECH_AOI222 U310 ( .A(n315), .B(n293), .C(n295), .D(n316), .E(n297), .F(
        n317), .Z(n314) );
  GTECH_NOT U311 ( .A(n318), .Z(N146) );
  GTECH_AOI222 U312 ( .A(n319), .B(n293), .C(n295), .D(n320), .E(n297), .F(
        n321), .Z(n318) );
  GTECH_NOT U313 ( .A(n322), .Z(N145) );
  GTECH_AOI222 U314 ( .A(n323), .B(n293), .C(n295), .D(n324), .E(n297), .F(
        n325), .Z(n322) );
  GTECH_NOT U315 ( .A(n326), .Z(N144) );
  GTECH_AOI222 U316 ( .A(n327), .B(n293), .C(n295), .D(n328), .E(n297), .F(
        n329), .Z(n326) );
  GTECH_NOT U317 ( .A(n330), .Z(N143) );
  GTECH_AOI222 U318 ( .A(n331), .B(n293), .C(n295), .D(n332), .E(n297), .F(
        n333), .Z(n330) );
  GTECH_NOT U319 ( .A(n334), .Z(N142) );
  GTECH_AOI222 U320 ( .A(n335), .B(n293), .C(n295), .D(n336), .E(n297), .F(
        n337), .Z(n334) );
  GTECH_NOT U321 ( .A(n338), .Z(N141) );
  GTECH_AOI222 U322 ( .A(n339), .B(n293), .C(n295), .D(n340), .E(n297), .F(
        n341), .Z(n338) );
  GTECH_NOT U323 ( .A(n342), .Z(N140) );
  GTECH_AOI222 U324 ( .A(n343), .B(n293), .C(n295), .D(n344), .E(n297), .F(
        n345), .Z(n342) );
  GTECH_NOT U325 ( .A(n346), .Z(N14) );
  GTECH_OR_NOT U326 ( .A(n305), .B(n287), .Z(n346) );
  GTECH_NOT U327 ( .A(n347), .Z(N139) );
  GTECH_AOI222 U328 ( .A(n348), .B(n293), .C(n295), .D(n349), .E(n297), .F(
        n350), .Z(n347) );
  GTECH_NOT U329 ( .A(n351), .Z(N138) );
  GTECH_AOI222 U330 ( .A(n352), .B(n293), .C(n295), .D(n353), .E(n297), .F(
        n354), .Z(n351) );
  GTECH_NOT U331 ( .A(n355), .Z(N137) );
  GTECH_AOI222 U332 ( .A(n356), .B(n293), .C(n295), .D(n357), .E(n297), .F(
        n358), .Z(n355) );
  GTECH_NOT U333 ( .A(n359), .Z(N136) );
  GTECH_AOI222 U334 ( .A(n293), .B(n272), .C(n295), .D(n274), .E(n297), .F(
        n276), .Z(n359) );
  GTECH_NOT U335 ( .A(n360), .Z(n276) );
  GTECH_XOR2 U336 ( .A(n361), .B(n362), .Z(n360) );
  GTECH_NOT U337 ( .A(n363), .Z(n362) );
  GTECH_NOT U338 ( .A(n364), .Z(n295) );
  GTECH_NOT U339 ( .A(n365), .Z(n272) );
  GTECH_XOR2 U340 ( .A(n361), .B(n366), .Z(n365) );
  GTECH_NOT U341 ( .A(n367), .Z(n366) );
  GTECH_XOR2 U342 ( .A(n274), .B(n254), .Z(n361) );
  GTECH_OAI21 U343 ( .A(n12), .B(n364), .C(n368), .Z(N135) );
  GTECH_OAI21 U344 ( .A(n297), .B(n293), .C(n280), .Z(n368) );
  GTECH_OAI21 U345 ( .A(n12), .B(n369), .C(n363), .Z(n280) );
  GTECH_NOT U346 ( .A(n253), .Z(n369) );
  GTECH_NOT U347 ( .A(n370), .Z(n293) );
  GTECH_OR3 U348 ( .A(n10), .B(n371), .C(n372), .Z(n370) );
  GTECH_NOT U349 ( .A(n373), .Z(n297) );
  GTECH_OR3 U350 ( .A(n28), .B(n374), .C(n372), .Z(n373) );
  GTECH_OR_NOT U351 ( .A(n372), .B(n375), .Z(n364) );
  GTECH_XOR2 U352 ( .A(n374), .B(n28), .Z(n375) );
  GTECH_AND2 U353 ( .A(N155), .B(n376), .Z(N134) );
  GTECH_NOT U354 ( .A(n13), .Z(n376) );
  GTECH_AND2 U355 ( .A(N155), .B(n377), .Z(N133) );
  GTECH_NOT U356 ( .A(n14), .Z(n377) );
  GTECH_AND2 U357 ( .A(N155), .B(n378), .Z(N132) );
  GTECH_NOT U358 ( .A(n15), .Z(n378) );
  GTECH_AND2 U359 ( .A(N155), .B(n379), .Z(N131) );
  GTECH_NOT U360 ( .A(n16), .Z(n379) );
  GTECH_AND2 U361 ( .A(N155), .B(n380), .Z(N130) );
  GTECH_NOT U362 ( .A(n17), .Z(n380) );
  GTECH_AND2 U363 ( .A(N155), .B(n381), .Z(N129) );
  GTECH_NOT U364 ( .A(n18), .Z(n381) );
  GTECH_AND2 U365 ( .A(N155), .B(n382), .Z(N128) );
  GTECH_NOT U366 ( .A(n19), .Z(n382) );
  GTECH_AND2 U367 ( .A(N155), .B(n383), .Z(N127) );
  GTECH_NOT U368 ( .A(n20), .Z(n383) );
  GTECH_AND2 U369 ( .A(N155), .B(n384), .Z(N126) );
  GTECH_NOT U370 ( .A(n21), .Z(n384) );
  GTECH_AND2 U371 ( .A(N155), .B(n385), .Z(N125) );
  GTECH_NOT U372 ( .A(n22), .Z(n385) );
  GTECH_AND2 U373 ( .A(N155), .B(n386), .Z(N124) );
  GTECH_NOT U374 ( .A(n23), .Z(n386) );
  GTECH_AND2 U375 ( .A(N155), .B(n387), .Z(N123) );
  GTECH_NOT U376 ( .A(n24), .Z(n387) );
  GTECH_AND2 U377 ( .A(N155), .B(n388), .Z(N122) );
  GTECH_NOT U378 ( .A(n25), .Z(n388) );
  GTECH_AND2 U379 ( .A(N155), .B(n389), .Z(N121) );
  GTECH_NOT U380 ( .A(n26), .Z(n389) );
  GTECH_AND2 U381 ( .A(N155), .B(n390), .Z(N120) );
  GTECH_NOT U382 ( .A(n27), .Z(n390) );
  GTECH_NOT U383 ( .A(n372), .Z(N155) );
  GTECH_NAND4 U384 ( .A(n8), .B(n7), .C(n9), .D(n391), .Z(n372) );
  GTECH_AND3 U385 ( .A(n299), .B(n305), .C(n6), .Z(n391) );
  GTECH_NOT U386 ( .A(n392), .Z(N116) );
  GTECH_AOI222 U387 ( .A(n273), .B(n296), .C(n275), .D(n298), .E(n294), .F(
        n271), .Z(n392) );
  GTECH_XOR2 U388 ( .A(n393), .B(n394), .Z(n294) );
  GTECH_ADD_ABC U389 ( .A(n31), .B(n268), .C(n395), .COUT(n394) );
  GTECH_XOR2 U390 ( .A(n396), .B(n393), .Z(n298) );
  GTECH_XOR2 U391 ( .A(A[16]), .B(n30), .Z(n393) );
  GTECH_OAI21 U392 ( .A(n397), .B(n31), .C(n398), .Z(n396) );
  GTECH_OAI21 U393 ( .A(n268), .B(n302), .C(n399), .Z(n398) );
  GTECH_NOT U394 ( .A(n30), .Z(n296) );
  GTECH_OR_NOT U395 ( .A(N41), .B(n283), .Z(N115) );
  GTECH_OR_NOT U396 ( .A(n281), .B(n299), .Z(N41) );
  GTECH_NOT U397 ( .A(Rst), .Z(n299) );
  GTECH_NOT U398 ( .A(n285), .Z(n281) );
  GTECH_OR_NOT U399 ( .A(Rst), .B(Ld), .Z(n285) );
  GTECH_NOT U400 ( .A(n400), .Z(N113) );
  GTECH_AOI222 U401 ( .A(n273), .B(n302), .C(n275), .D(n303), .E(n301), .F(
        n271), .Z(n400) );
  GTECH_XOR2 U402 ( .A(n401), .B(n395), .Z(n301) );
  GTECH_ADD_ABC U403 ( .A(n32), .B(n267), .C(n402), .COUT(n395) );
  GTECH_NOT U404 ( .A(n403), .Z(n303) );
  GTECH_XOR2 U405 ( .A(n401), .B(n404), .Z(n403) );
  GTECH_NOT U406 ( .A(n399), .Z(n404) );
  GTECH_OAI21 U407 ( .A(n32), .B(n405), .C(n406), .Z(n399) );
  GTECH_OAI21 U408 ( .A(n267), .B(n308), .C(n407), .Z(n406) );
  GTECH_XOR2 U409 ( .A(n397), .B(n31), .Z(n401) );
  GTECH_NOT U410 ( .A(n268), .Z(n397) );
  GTECH_NOT U411 ( .A(n31), .Z(n302) );
  GTECH_NOT U412 ( .A(n408), .Z(N112) );
  GTECH_AOI222 U413 ( .A(n273), .B(n308), .C(n275), .D(n309), .E(n307), .F(
        n271), .Z(n408) );
  GTECH_XOR2 U414 ( .A(n409), .B(n402), .Z(n307) );
  GTECH_ADD_ABC U415 ( .A(n33), .B(n266), .C(n410), .COUT(n402) );
  GTECH_NOT U416 ( .A(n411), .Z(n309) );
  GTECH_XOR2 U417 ( .A(n409), .B(n412), .Z(n411) );
  GTECH_NOT U418 ( .A(n407), .Z(n412) );
  GTECH_OAI21 U419 ( .A(n33), .B(n413), .C(n414), .Z(n407) );
  GTECH_OAI21 U420 ( .A(n266), .B(n312), .C(n415), .Z(n414) );
  GTECH_XOR2 U421 ( .A(n405), .B(n32), .Z(n409) );
  GTECH_NOT U422 ( .A(n267), .Z(n405) );
  GTECH_NOT U423 ( .A(n32), .Z(n308) );
  GTECH_NOT U424 ( .A(n416), .Z(N111) );
  GTECH_AOI222 U425 ( .A(n273), .B(n312), .C(n275), .D(n313), .E(n311), .F(
        n271), .Z(n416) );
  GTECH_XOR2 U426 ( .A(n417), .B(n410), .Z(n311) );
  GTECH_ADD_ABC U427 ( .A(n34), .B(n265), .C(n418), .COUT(n410) );
  GTECH_NOT U428 ( .A(n419), .Z(n313) );
  GTECH_XOR2 U429 ( .A(n417), .B(n420), .Z(n419) );
  GTECH_NOT U430 ( .A(n415), .Z(n420) );
  GTECH_OAI21 U431 ( .A(n34), .B(n421), .C(n422), .Z(n415) );
  GTECH_OAI21 U432 ( .A(n265), .B(n316), .C(n423), .Z(n422) );
  GTECH_XOR2 U433 ( .A(n413), .B(n33), .Z(n417) );
  GTECH_NOT U434 ( .A(n266), .Z(n413) );
  GTECH_NOT U435 ( .A(n33), .Z(n312) );
  GTECH_NOT U436 ( .A(n424), .Z(N110) );
  GTECH_AOI222 U437 ( .A(n273), .B(n316), .C(n275), .D(n317), .E(n315), .F(
        n271), .Z(n424) );
  GTECH_XOR2 U438 ( .A(n425), .B(n418), .Z(n315) );
  GTECH_ADD_ABC U439 ( .A(n35), .B(n264), .C(n426), .COUT(n418) );
  GTECH_NOT U440 ( .A(n427), .Z(n317) );
  GTECH_XOR2 U441 ( .A(n425), .B(n428), .Z(n427) );
  GTECH_NOT U442 ( .A(n423), .Z(n428) );
  GTECH_OAI21 U443 ( .A(n35), .B(n429), .C(n430), .Z(n423) );
  GTECH_OAI21 U444 ( .A(n264), .B(n320), .C(n431), .Z(n430) );
  GTECH_XOR2 U445 ( .A(n421), .B(n34), .Z(n425) );
  GTECH_NOT U446 ( .A(n265), .Z(n421) );
  GTECH_NOT U447 ( .A(n34), .Z(n316) );
  GTECH_NOT U448 ( .A(n432), .Z(N109) );
  GTECH_AOI222 U449 ( .A(n273), .B(n320), .C(n275), .D(n321), .E(n319), .F(
        n271), .Z(n432) );
  GTECH_XOR2 U450 ( .A(n433), .B(n426), .Z(n319) );
  GTECH_ADD_ABC U451 ( .A(n36), .B(n263), .C(n434), .COUT(n426) );
  GTECH_NOT U452 ( .A(n435), .Z(n321) );
  GTECH_XOR2 U453 ( .A(n433), .B(n436), .Z(n435) );
  GTECH_NOT U454 ( .A(n431), .Z(n436) );
  GTECH_OAI21 U455 ( .A(n36), .B(n437), .C(n438), .Z(n431) );
  GTECH_OAI21 U456 ( .A(n263), .B(n324), .C(n439), .Z(n438) );
  GTECH_XOR2 U457 ( .A(n429), .B(n35), .Z(n433) );
  GTECH_NOT U458 ( .A(n264), .Z(n429) );
  GTECH_NOT U459 ( .A(n35), .Z(n320) );
  GTECH_NOT U460 ( .A(n440), .Z(N108) );
  GTECH_AOI222 U461 ( .A(n273), .B(n324), .C(n275), .D(n325), .E(n323), .F(
        n271), .Z(n440) );
  GTECH_XOR2 U462 ( .A(n441), .B(n434), .Z(n323) );
  GTECH_ADD_ABC U463 ( .A(n37), .B(n262), .C(n442), .COUT(n434) );
  GTECH_NOT U464 ( .A(n443), .Z(n325) );
  GTECH_XOR2 U465 ( .A(n441), .B(n444), .Z(n443) );
  GTECH_NOT U466 ( .A(n439), .Z(n444) );
  GTECH_OAI21 U467 ( .A(n37), .B(n445), .C(n446), .Z(n439) );
  GTECH_OAI21 U468 ( .A(n262), .B(n328), .C(n447), .Z(n446) );
  GTECH_XOR2 U469 ( .A(n437), .B(n36), .Z(n441) );
  GTECH_NOT U470 ( .A(n263), .Z(n437) );
  GTECH_NOT U471 ( .A(n36), .Z(n324) );
  GTECH_NOT U472 ( .A(n448), .Z(N107) );
  GTECH_AOI222 U473 ( .A(n273), .B(n328), .C(n275), .D(n329), .E(n327), .F(
        n271), .Z(n448) );
  GTECH_XOR2 U474 ( .A(n449), .B(n442), .Z(n327) );
  GTECH_ADD_ABC U475 ( .A(n38), .B(n261), .C(n450), .COUT(n442) );
  GTECH_NOT U476 ( .A(n451), .Z(n329) );
  GTECH_XOR2 U477 ( .A(n449), .B(n452), .Z(n451) );
  GTECH_NOT U478 ( .A(n447), .Z(n452) );
  GTECH_OAI21 U479 ( .A(n38), .B(n453), .C(n454), .Z(n447) );
  GTECH_OAI21 U480 ( .A(n261), .B(n332), .C(n455), .Z(n454) );
  GTECH_XOR2 U481 ( .A(n445), .B(n37), .Z(n449) );
  GTECH_NOT U482 ( .A(n262), .Z(n445) );
  GTECH_NOT U483 ( .A(n37), .Z(n328) );
  GTECH_NOT U484 ( .A(n456), .Z(N106) );
  GTECH_AOI222 U485 ( .A(n273), .B(n332), .C(n275), .D(n333), .E(n331), .F(
        n271), .Z(n456) );
  GTECH_XOR2 U486 ( .A(n457), .B(n450), .Z(n331) );
  GTECH_ADD_ABC U487 ( .A(n39), .B(n260), .C(n458), .COUT(n450) );
  GTECH_NOT U488 ( .A(n459), .Z(n333) );
  GTECH_XOR2 U489 ( .A(n457), .B(n460), .Z(n459) );
  GTECH_NOT U490 ( .A(n455), .Z(n460) );
  GTECH_OAI21 U491 ( .A(n39), .B(n461), .C(n462), .Z(n455) );
  GTECH_OAI21 U492 ( .A(n260), .B(n336), .C(n463), .Z(n462) );
  GTECH_XOR2 U493 ( .A(n453), .B(n38), .Z(n457) );
  GTECH_NOT U494 ( .A(n261), .Z(n453) );
  GTECH_NOT U495 ( .A(n38), .Z(n332) );
  GTECH_NOT U496 ( .A(n464), .Z(N105) );
  GTECH_AOI222 U497 ( .A(n273), .B(n336), .C(n275), .D(n337), .E(n335), .F(
        n271), .Z(n464) );
  GTECH_XOR2 U498 ( .A(n465), .B(n458), .Z(n335) );
  GTECH_ADD_ABC U499 ( .A(n40), .B(n259), .C(n466), .COUT(n458) );
  GTECH_NOT U500 ( .A(n467), .Z(n337) );
  GTECH_XOR2 U501 ( .A(n465), .B(n468), .Z(n467) );
  GTECH_NOT U502 ( .A(n463), .Z(n468) );
  GTECH_OAI21 U503 ( .A(n40), .B(n469), .C(n470), .Z(n463) );
  GTECH_OAI21 U504 ( .A(n259), .B(n340), .C(n471), .Z(n470) );
  GTECH_XOR2 U505 ( .A(n461), .B(n39), .Z(n465) );
  GTECH_NOT U506 ( .A(n260), .Z(n461) );
  GTECH_NOT U507 ( .A(n39), .Z(n336) );
  GTECH_NOT U508 ( .A(n472), .Z(N104) );
  GTECH_AOI222 U509 ( .A(n273), .B(n340), .C(n275), .D(n341), .E(n339), .F(
        n271), .Z(n472) );
  GTECH_XOR2 U510 ( .A(n473), .B(n466), .Z(n339) );
  GTECH_ADD_ABC U511 ( .A(n41), .B(n258), .C(n474), .COUT(n466) );
  GTECH_NOT U512 ( .A(n475), .Z(n341) );
  GTECH_XOR2 U513 ( .A(n473), .B(n476), .Z(n475) );
  GTECH_NOT U514 ( .A(n471), .Z(n476) );
  GTECH_OAI21 U515 ( .A(n41), .B(n477), .C(n478), .Z(n471) );
  GTECH_OAI21 U516 ( .A(n258), .B(n344), .C(n479), .Z(n478) );
  GTECH_XOR2 U517 ( .A(n469), .B(n40), .Z(n473) );
  GTECH_NOT U518 ( .A(n259), .Z(n469) );
  GTECH_NOT U519 ( .A(n40), .Z(n340) );
  GTECH_NOT U520 ( .A(n480), .Z(N103) );
  GTECH_AOI222 U521 ( .A(n273), .B(n344), .C(n275), .D(n345), .E(n343), .F(
        n271), .Z(n480) );
  GTECH_XOR2 U522 ( .A(n481), .B(n474), .Z(n343) );
  GTECH_ADD_ABC U523 ( .A(n42), .B(n257), .C(n482), .COUT(n474) );
  GTECH_NOT U524 ( .A(n483), .Z(n345) );
  GTECH_XOR2 U525 ( .A(n481), .B(n484), .Z(n483) );
  GTECH_NOT U526 ( .A(n479), .Z(n484) );
  GTECH_OAI21 U527 ( .A(n42), .B(n485), .C(n486), .Z(n479) );
  GTECH_OAI21 U528 ( .A(n257), .B(n349), .C(n487), .Z(n486) );
  GTECH_XOR2 U529 ( .A(n477), .B(n41), .Z(n481) );
  GTECH_NOT U530 ( .A(n258), .Z(n477) );
  GTECH_NOT U531 ( .A(n41), .Z(n344) );
  GTECH_NOT U532 ( .A(n488), .Z(N102) );
  GTECH_AOI222 U533 ( .A(n273), .B(n349), .C(n275), .D(n350), .E(n348), .F(
        n271), .Z(n488) );
  GTECH_XOR2 U534 ( .A(n489), .B(n482), .Z(n348) );
  GTECH_ADD_ABC U535 ( .A(n43), .B(n256), .C(n490), .COUT(n482) );
  GTECH_NOT U536 ( .A(n491), .Z(n350) );
  GTECH_XOR2 U537 ( .A(n489), .B(n492), .Z(n491) );
  GTECH_NOT U538 ( .A(n487), .Z(n492) );
  GTECH_OAI21 U539 ( .A(n43), .B(n493), .C(n494), .Z(n487) );
  GTECH_OAI21 U540 ( .A(n256), .B(n353), .C(n495), .Z(n494) );
  GTECH_XOR2 U541 ( .A(n485), .B(n42), .Z(n489) );
  GTECH_NOT U542 ( .A(n257), .Z(n485) );
  GTECH_NOT U543 ( .A(n42), .Z(n349) );
  GTECH_NOT U544 ( .A(n496), .Z(N101) );
  GTECH_AOI222 U545 ( .A(n273), .B(n353), .C(n275), .D(n354), .E(n352), .F(
        n271), .Z(n496) );
  GTECH_XOR2 U546 ( .A(n497), .B(n490), .Z(n352) );
  GTECH_ADD_ABC U547 ( .A(n29), .B(n255), .C(n498), .COUT(n490) );
  GTECH_NOT U548 ( .A(n499), .Z(n354) );
  GTECH_XOR2 U549 ( .A(n497), .B(n500), .Z(n499) );
  GTECH_NOT U550 ( .A(n495), .Z(n500) );
  GTECH_OAI21 U551 ( .A(n29), .B(n501), .C(n502), .Z(n495) );
  GTECH_OAI21 U552 ( .A(n255), .B(n357), .C(n503), .Z(n502) );
  GTECH_XOR2 U553 ( .A(n493), .B(n43), .Z(n497) );
  GTECH_NOT U554 ( .A(n256), .Z(n493) );
  GTECH_NOT U555 ( .A(n43), .Z(n353) );
  GTECH_NOT U556 ( .A(n504), .Z(N100) );
  GTECH_AOI222 U557 ( .A(n356), .B(n271), .C(n273), .D(n357), .E(n275), .F(
        n358), .Z(n504) );
  GTECH_NOT U558 ( .A(n505), .Z(n358) );
  GTECH_XOR2 U559 ( .A(n506), .B(n507), .Z(n505) );
  GTECH_NOT U560 ( .A(n503), .Z(n507) );
  GTECH_OAI21 U561 ( .A(n11), .B(n508), .C(n509), .Z(n503) );
  GTECH_OAI21 U562 ( .A(n254), .B(n274), .C(n363), .Z(n509) );
  GTECH_OR_NOT U563 ( .A(n253), .B(n12), .Z(n363) );
  GTECH_NOT U564 ( .A(n11), .Z(n274) );
  GTECH_NOT U565 ( .A(n254), .Z(n508) );
  GTECH_NOT U566 ( .A(n510), .Z(n275) );
  GTECH_OR_NOT U567 ( .A(n374), .B(N82), .Z(n510) );
  GTECH_NOT U568 ( .A(n511), .Z(N82) );
  GTECH_NOT U569 ( .A(n10), .Z(n374) );
  GTECH_NOT U570 ( .A(n29), .Z(n357) );
  GTECH_NOT U571 ( .A(n512), .Z(n273) );
  GTECH_MUX2 U572 ( .A(n511), .B(n513), .S(n10), .Z(n512) );
  GTECH_OR_NOT U573 ( .A(n283), .B(n28), .Z(n513) );
  GTECH_OR_NOT U574 ( .A(n28), .B(n287), .Z(n511) );
  GTECH_NOT U575 ( .A(n283), .Z(n287) );
  GTECH_NOT U576 ( .A(n282), .Z(n271) );
  GTECH_OR3 U577 ( .A(n10), .B(n283), .C(n371), .Z(n282) );
  GTECH_NOT U578 ( .A(n28), .Z(n371) );
  GTECH_OR3 U579 ( .A(Ld), .B(Rst), .C(n514), .Z(n283) );
  GTECH_AND_NOT U580 ( .A(n9), .B(n286), .Z(n514) );
  GTECH_OR_NOT U581 ( .A(n289), .B(n8), .Z(n286) );
  GTECH_OR_NOT U582 ( .A(n291), .B(n7), .Z(n289) );
  GTECH_OR_NOT U583 ( .A(n305), .B(n6), .Z(n291) );
  GTECH_NOT U584 ( .A(n252), .Z(n305) );
  GTECH_XOR2 U585 ( .A(n506), .B(n498), .Z(n356) );
  GTECH_ADD_ABC U586 ( .A(n254), .B(n11), .C(n367), .COUT(n498) );
  GTECH_OR_NOT U587 ( .A(n253), .B(n278), .Z(n367) );
  GTECH_NOT U588 ( .A(n12), .Z(n278) );
  GTECH_XOR2 U589 ( .A(n501), .B(n29), .Z(n506) );
  GTECH_NOT U590 ( .A(n255), .Z(n501) );
endmodule

