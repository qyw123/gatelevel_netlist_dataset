
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n113, n114, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK2S Cntr_reg_0_ ( .J(n114), .K(n114), .TI(N14), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[0]), .QN(n338) );
  GTECH_FJK2S Cntr_reg_1_ ( .J(n114), .K(n114), .TI(N15), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK2S Cntr_reg_2_ ( .J(n114), .K(n114), .TI(N16), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK2S Cntr_reg_3_ ( .J(n114), .K(n114), .TI(N17), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK2S Cntr_reg_4_ ( .J(n114), .K(n114), .TI(N19), .TE(N18), .CP(clk), 
        .CD(n113), .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK2S A_reg_16_ ( .J(n114), .K(n114), .TI(N42), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[16]), .QN(n355) );
  GTECH_FJK2S A_reg_15_ ( .J(n114), .K(n114), .TI(N42), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[15]), .QN(n354) );
  GTECH_FJK2S A_reg_14_ ( .J(n114), .K(n114), .TI(N39), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[14]), .QN(n353) );
  GTECH_FJK2S A_reg_13_ ( .J(n114), .K(n114), .TI(N38), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[13]), .QN(n352) );
  GTECH_FJK2S A_reg_12_ ( .J(n114), .K(n114), .TI(N37), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[12]), .QN(n351) );
  GTECH_FJK2S A_reg_11_ ( .J(n114), .K(n114), .TI(N36), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[11]), .QN(n350) );
  GTECH_FJK2S A_reg_10_ ( .J(n114), .K(n114), .TI(N35), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[10]), .QN(n349) );
  GTECH_FJK2S A_reg_9_ ( .J(n114), .K(n114), .TI(N34), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[9]), .QN(n348) );
  GTECH_FJK2S A_reg_8_ ( .J(n114), .K(n114), .TI(N33), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[8]), .QN(n347) );
  GTECH_FJK2S A_reg_7_ ( .J(n114), .K(n114), .TI(N32), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[7]), .QN(n346) );
  GTECH_FJK2S A_reg_6_ ( .J(n114), .K(n114), .TI(N31), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[6]), .QN(n345) );
  GTECH_FJK2S A_reg_5_ ( .J(n114), .K(n114), .TI(N30), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[5]), .QN(n344) );
  GTECH_FJK2S A_reg_4_ ( .J(n114), .K(n114), .TI(N29), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[4]), .QN(n343) );
  GTECH_FJK2S A_reg_3_ ( .J(n114), .K(n114), .TI(N28), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[3]), .QN(n342) );
  GTECH_FJK2S A_reg_2_ ( .J(n114), .K(n114), .TI(N27), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[2]), .QN(n341) );
  GTECH_FJK2S A_reg_1_ ( .J(n114), .K(n114), .TI(N26), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[1]), .QN(n340) );
  GTECH_FJK2S A_reg_0_ ( .J(n114), .K(n114), .TI(N25), .TE(N41), .CP(clk), 
        .CD(n113), .Q(A[0]), .QN(n339) );
  GTECH_FJK2S Prod_reg_0_ ( .J(n114), .K(n114), .TI(N82), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[0]), .QN(n10) );
  GTECH_FJK2S Prod_reg_18_ ( .J(n114), .K(n114), .TI(N100), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK2S Prod_reg_17_ ( .J(n114), .K(n114), .TI(N99), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[17]), .QN(n12) );
  GTECH_FJK2S Prod_reg_16_ ( .J(n114), .K(n114), .TI(N98), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[16]), .QN(n13) );
  GTECH_FJK2S Prod_reg_15_ ( .J(n114), .K(n114), .TI(N97), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[15]), .QN(n14) );
  GTECH_FJK2S Prod_reg_14_ ( .J(n114), .K(n114), .TI(N96), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[14]), .QN(n15) );
  GTECH_FJK2S Prod_reg_13_ ( .J(n114), .K(n114), .TI(N95), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[13]), .QN(n16) );
  GTECH_FJK2S Prod_reg_12_ ( .J(n114), .K(n114), .TI(N94), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[12]), .QN(n17) );
  GTECH_FJK2S Prod_reg_11_ ( .J(n114), .K(n114), .TI(N93), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[11]), .QN(n18) );
  GTECH_FJK2S Prod_reg_10_ ( .J(n114), .K(n114), .TI(N92), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[10]), .QN(n19) );
  GTECH_FJK2S Prod_reg_9_ ( .J(n114), .K(n114), .TI(N91), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[9]), .QN(n20) );
  GTECH_FJK2S Prod_reg_8_ ( .J(n114), .K(n114), .TI(N90), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[8]), .QN(n21) );
  GTECH_FJK2S Prod_reg_7_ ( .J(n114), .K(n114), .TI(N89), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[7]), .QN(n22) );
  GTECH_FJK2S Prod_reg_6_ ( .J(n114), .K(n114), .TI(N88), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[6]), .QN(n23) );
  GTECH_FJK2S Prod_reg_5_ ( .J(n114), .K(n114), .TI(N87), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[5]), .QN(n24) );
  GTECH_FJK2S Prod_reg_4_ ( .J(n114), .K(n114), .TI(N86), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[4]), .QN(n25) );
  GTECH_FJK2S Prod_reg_3_ ( .J(n114), .K(n114), .TI(N85), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[3]), .QN(n26) );
  GTECH_FJK2S Prod_reg_2_ ( .J(n114), .K(n114), .TI(N84), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[2]), .QN(n27) );
  GTECH_FJK2S Prod_reg_1_ ( .J(n114), .K(n114), .TI(N83), .TE(N115), .CP(clk), 
        .CD(n113), .Q(Prod[1]), .QN(n28) );
  GTECH_FJK2S Prod_reg_19_ ( .J(n114), .K(n114), .TI(N101), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK2S Prod_reg_33_ ( .J(n114), .K(n114), .TI(N116), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK2S Prod_reg_32_ ( .J(n114), .K(n114), .TI(N116), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK2S Prod_reg_31_ ( .J(n114), .K(n114), .TI(N113), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK2S Prod_reg_30_ ( .J(n114), .K(n114), .TI(N112), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK2S Prod_reg_29_ ( .J(n114), .K(n114), .TI(N111), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK2S Prod_reg_28_ ( .J(n114), .K(n114), .TI(N110), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK2S Prod_reg_27_ ( .J(n114), .K(n114), .TI(N109), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK2S Prod_reg_26_ ( .J(n114), .K(n114), .TI(N108), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK2S Prod_reg_25_ ( .J(n114), .K(n114), .TI(N107), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK2S Prod_reg_24_ ( .J(n114), .K(n114), .TI(N106), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK2S Prod_reg_23_ ( .J(n114), .K(n114), .TI(N105), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK2S Prod_reg_22_ ( .J(n114), .K(n114), .TI(N104), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK2S Prod_reg_21_ ( .J(n114), .K(n114), .TI(N103), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK2S Prod_reg_20_ ( .J(n114), .K(n114), .TI(N102), .TE(N115), .CP(clk), .CD(n113), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK2S P_reg_31_ ( .J(n114), .K(n114), .TI(N152), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[31]) );
  GTECH_FJK2S P_reg_30_ ( .J(n114), .K(n114), .TI(N150), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[30]) );
  GTECH_FJK2S P_reg_29_ ( .J(n114), .K(n114), .TI(N149), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[29]) );
  GTECH_FJK2S P_reg_28_ ( .J(n114), .K(n114), .TI(N148), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[28]) );
  GTECH_FJK2S P_reg_27_ ( .J(n114), .K(n114), .TI(N147), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[27]) );
  GTECH_FJK2S P_reg_26_ ( .J(n114), .K(n114), .TI(N146), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[26]) );
  GTECH_FJK2S P_reg_25_ ( .J(n114), .K(n114), .TI(N145), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[25]) );
  GTECH_FJK2S P_reg_24_ ( .J(n114), .K(n114), .TI(N144), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[24]) );
  GTECH_FJK2S P_reg_23_ ( .J(n114), .K(n114), .TI(N143), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[23]) );
  GTECH_FJK2S P_reg_22_ ( .J(n114), .K(n114), .TI(N142), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[22]) );
  GTECH_FJK2S P_reg_21_ ( .J(n114), .K(n114), .TI(N141), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[21]) );
  GTECH_FJK2S P_reg_20_ ( .J(n114), .K(n114), .TI(N140), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[20]) );
  GTECH_FJK2S P_reg_19_ ( .J(n114), .K(n114), .TI(N139), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[19]) );
  GTECH_FJK2S P_reg_18_ ( .J(n114), .K(n114), .TI(N138), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[18]) );
  GTECH_FJK2S P_reg_17_ ( .J(n114), .K(n114), .TI(N137), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[17]) );
  GTECH_FJK2S P_reg_16_ ( .J(n114), .K(n114), .TI(N136), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[16]) );
  GTECH_FJK2S P_reg_15_ ( .J(n114), .K(n114), .TI(N135), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[15]) );
  GTECH_FJK2S P_reg_14_ ( .J(n114), .K(n114), .TI(N134), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[14]) );
  GTECH_FJK2S P_reg_13_ ( .J(n114), .K(n114), .TI(N133), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[13]) );
  GTECH_FJK2S P_reg_12_ ( .J(n114), .K(n114), .TI(N132), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[12]) );
  GTECH_FJK2S P_reg_11_ ( .J(n114), .K(n114), .TI(N131), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[11]) );
  GTECH_FJK2S P_reg_10_ ( .J(n114), .K(n114), .TI(N130), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[10]) );
  GTECH_FJK2S P_reg_9_ ( .J(n114), .K(n114), .TI(N129), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[9]) );
  GTECH_FJK2S P_reg_8_ ( .J(n114), .K(n114), .TI(N128), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[8]) );
  GTECH_FJK2S P_reg_7_ ( .J(n114), .K(n114), .TI(N127), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[7]) );
  GTECH_FJK2S P_reg_6_ ( .J(n114), .K(n114), .TI(N126), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[6]) );
  GTECH_FJK2S P_reg_5_ ( .J(n114), .K(n114), .TI(N125), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[5]) );
  GTECH_FJK2S P_reg_4_ ( .J(n114), .K(n114), .TI(N124), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[4]) );
  GTECH_FJK2S P_reg_3_ ( .J(n114), .K(n114), .TI(N123), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[3]) );
  GTECH_FJK2S P_reg_2_ ( .J(n114), .K(n114), .TI(N122), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[2]) );
  GTECH_FJK2S P_reg_1_ ( .J(n114), .K(n114), .TI(N121), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[1]) );
  GTECH_FJK2S P_reg_0_ ( .J(n114), .K(n114), .TI(N120), .TE(N151), .CP(clk), 
        .CD(n113), .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U340 ( .Z(n114) );
  GTECH_ONE U341 ( .Z(n113) );
  GTECH_NOT U342 ( .A(n356), .Z(N99) );
  GTECH_AOI222 U343 ( .A(n357), .B(n358), .C(n359), .D(n360), .E(n361), .F(
        n362), .Z(n356) );
  GTECH_NOT U344 ( .A(n363), .Z(N98) );
  GTECH_AOI222 U345 ( .A(n359), .B(n364), .C(n365), .D(n366), .E(R[15]), .F(
        n367), .Z(n363) );
  GTECH_NAND2 U346 ( .A(n368), .B(n369), .Z(n365) );
  GTECH_OAI2N2 U347 ( .A(n13), .B(n370), .C(R[14]), .D(n367), .Z(N97) );
  GTECH_OAI2N2 U348 ( .A(n14), .B(n370), .C(R[13]), .D(n367), .Z(N96) );
  GTECH_OAI2N2 U349 ( .A(n15), .B(n370), .C(R[12]), .D(n367), .Z(N95) );
  GTECH_OAI2N2 U350 ( .A(n16), .B(n370), .C(R[11]), .D(n367), .Z(N94) );
  GTECH_OAI2N2 U351 ( .A(n17), .B(n370), .C(R[10]), .D(n367), .Z(N93) );
  GTECH_OAI2N2 U352 ( .A(n18), .B(n370), .C(R[9]), .D(n367), .Z(N92) );
  GTECH_OAI2N2 U353 ( .A(n19), .B(n370), .C(R[8]), .D(n367), .Z(N91) );
  GTECH_OAI2N2 U354 ( .A(n20), .B(n370), .C(R[7]), .D(n367), .Z(N90) );
  GTECH_OAI2N2 U355 ( .A(n21), .B(n370), .C(R[6]), .D(n367), .Z(N89) );
  GTECH_OAI2N2 U356 ( .A(n22), .B(n370), .C(R[5]), .D(n367), .Z(N88) );
  GTECH_OAI2N2 U357 ( .A(n23), .B(n370), .C(R[4]), .D(n367), .Z(N87) );
  GTECH_OAI2N2 U358 ( .A(n24), .B(n370), .C(R[3]), .D(n367), .Z(N86) );
  GTECH_OAI2N2 U359 ( .A(n25), .B(n370), .C(R[2]), .D(n367), .Z(N85) );
  GTECH_OAI2N2 U360 ( .A(n26), .B(n370), .C(R[1]), .D(n367), .Z(N84) );
  GTECH_OAI2N2 U361 ( .A(n27), .B(n370), .C(R[0]), .D(n367), .Z(N83) );
  GTECH_AND2 U362 ( .A(M[15]), .B(n367), .Z(N42) );
  GTECH_AND2 U363 ( .A(M[14]), .B(n367), .Z(N39) );
  GTECH_AND2 U364 ( .A(M[13]), .B(n367), .Z(N38) );
  GTECH_AND2 U365 ( .A(M[12]), .B(n367), .Z(N37) );
  GTECH_AND2 U366 ( .A(M[11]), .B(n367), .Z(N36) );
  GTECH_AND2 U367 ( .A(M[10]), .B(n367), .Z(N35) );
  GTECH_AND2 U368 ( .A(M[9]), .B(n367), .Z(N34) );
  GTECH_AND2 U369 ( .A(M[8]), .B(n367), .Z(N33) );
  GTECH_AND2 U370 ( .A(M[7]), .B(n367), .Z(N32) );
  GTECH_AND2 U371 ( .A(M[6]), .B(n367), .Z(N31) );
  GTECH_AND2 U372 ( .A(M[5]), .B(n367), .Z(N30) );
  GTECH_AND2 U373 ( .A(M[4]), .B(n367), .Z(N29) );
  GTECH_AND2 U374 ( .A(M[3]), .B(n367), .Z(N28) );
  GTECH_AND2 U375 ( .A(M[2]), .B(n367), .Z(N27) );
  GTECH_AND2 U376 ( .A(M[1]), .B(n367), .Z(N26) );
  GTECH_AND2 U377 ( .A(M[0]), .B(n367), .Z(N25) );
  GTECH_NOT U378 ( .A(n371), .Z(n367) );
  GTECH_NAND2 U379 ( .A(n371), .B(n372), .Z(N19) );
  GTECH_NAND3 U380 ( .A(n373), .B(n374), .C(n375), .Z(n372) );
  GTECH_NAND3 U381 ( .A(n376), .B(n377), .C(n370), .Z(N18) );
  GTECH_AND2 U382 ( .A(n375), .B(n378), .Z(N17) );
  GTECH_OAI21 U383 ( .A(n8), .B(n379), .C(n373), .Z(n378) );
  GTECH_AND2 U384 ( .A(n375), .B(n380), .Z(N16) );
  GTECH_OAI21 U385 ( .A(n7), .B(n381), .C(n382), .Z(n380) );
  GTECH_NOT U386 ( .A(n383), .Z(N152) );
  GTECH_AOI222 U387 ( .A(n384), .B(n385), .C(n386), .D(n387), .E(n388), .F(
        n389), .Z(n383) );
  GTECH_NAND2 U388 ( .A(n377), .B(n390), .Z(N151) );
  GTECH_NOT U389 ( .A(n391), .Z(N150) );
  GTECH_AOI222 U390 ( .A(n392), .B(n384), .C(n386), .D(n393), .E(n388), .F(
        n394), .Z(n391) );
  GTECH_OAI21 U391 ( .A(n395), .B(n396), .C(n397), .Z(N15) );
  GTECH_NAND3 U392 ( .A(n375), .B(n398), .C(n395), .Z(n397) );
  GTECH_NOT U393 ( .A(n6), .Z(n395) );
  GTECH_NOT U394 ( .A(n399), .Z(N149) );
  GTECH_AOI222 U395 ( .A(n400), .B(n384), .C(n386), .D(n401), .E(n388), .F(
        n402), .Z(n399) );
  GTECH_NOT U396 ( .A(n403), .Z(N148) );
  GTECH_AOI222 U397 ( .A(n404), .B(n384), .C(n386), .D(n405), .E(n388), .F(
        n406), .Z(n403) );
  GTECH_NOT U398 ( .A(n407), .Z(N147) );
  GTECH_AOI222 U399 ( .A(n408), .B(n384), .C(n386), .D(n409), .E(n388), .F(
        n410), .Z(n407) );
  GTECH_NOT U400 ( .A(n411), .Z(N146) );
  GTECH_AOI222 U401 ( .A(n412), .B(n384), .C(n386), .D(n413), .E(n388), .F(
        n414), .Z(n411) );
  GTECH_NOT U402 ( .A(n415), .Z(N145) );
  GTECH_AOI222 U403 ( .A(n416), .B(n384), .C(n386), .D(n417), .E(n388), .F(
        n418), .Z(n415) );
  GTECH_NOT U404 ( .A(n419), .Z(N144) );
  GTECH_AOI222 U405 ( .A(n420), .B(n384), .C(n386), .D(n421), .E(n388), .F(
        n422), .Z(n419) );
  GTECH_NOT U406 ( .A(n423), .Z(N143) );
  GTECH_AOI222 U407 ( .A(n424), .B(n384), .C(n386), .D(n425), .E(n388), .F(
        n426), .Z(n423) );
  GTECH_NOT U408 ( .A(n427), .Z(N142) );
  GTECH_AOI222 U409 ( .A(n428), .B(n384), .C(n386), .D(n429), .E(n388), .F(
        n430), .Z(n427) );
  GTECH_NOT U410 ( .A(n431), .Z(N141) );
  GTECH_AOI222 U411 ( .A(n432), .B(n384), .C(n386), .D(n433), .E(n388), .F(
        n434), .Z(n431) );
  GTECH_NOT U412 ( .A(n435), .Z(N140) );
  GTECH_AOI222 U413 ( .A(n436), .B(n384), .C(n386), .D(n437), .E(n388), .F(
        n438), .Z(n435) );
  GTECH_NOT U414 ( .A(n396), .Z(N14) );
  GTECH_NAND2 U415 ( .A(n375), .B(n338), .Z(n396) );
  GTECH_NOT U416 ( .A(n439), .Z(N139) );
  GTECH_AOI222 U417 ( .A(n440), .B(n384), .C(n386), .D(n441), .E(n388), .F(
        n442), .Z(n439) );
  GTECH_NOT U418 ( .A(n443), .Z(N138) );
  GTECH_AOI222 U419 ( .A(n444), .B(n384), .C(n386), .D(n445), .E(n388), .F(
        n446), .Z(n443) );
  GTECH_NOT U420 ( .A(n447), .Z(N137) );
  GTECH_AOI222 U421 ( .A(n448), .B(n384), .C(n386), .D(n449), .E(n388), .F(
        n450), .Z(n447) );
  GTECH_NOT U422 ( .A(n451), .Z(N136) );
  GTECH_AOI222 U423 ( .A(n384), .B(n358), .C(n386), .D(n360), .E(n388), .F(
        n362), .Z(n451) );
  GTECH_NOT U424 ( .A(n452), .Z(n362) );
  GTECH_XOR2 U425 ( .A(n453), .B(n454), .Z(n452) );
  GTECH_NOT U426 ( .A(n455), .Z(n454) );
  GTECH_NOT U427 ( .A(n456), .Z(n386) );
  GTECH_NOT U428 ( .A(n457), .Z(n358) );
  GTECH_XOR2 U429 ( .A(n453), .B(n458), .Z(n457) );
  GTECH_NOT U430 ( .A(n459), .Z(n458) );
  GTECH_XOR2 U431 ( .A(n360), .B(n340), .Z(n453) );
  GTECH_OAI21 U432 ( .A(n12), .B(n456), .C(n460), .Z(N135) );
  GTECH_OAI21 U433 ( .A(n388), .B(n384), .C(n366), .Z(n460) );
  GTECH_OAI21 U434 ( .A(n12), .B(n461), .C(n455), .Z(n366) );
  GTECH_NOT U435 ( .A(n462), .Z(n384) );
  GTECH_NAND3 U436 ( .A(n28), .B(n463), .C(N155), .Z(n462) );
  GTECH_NOT U437 ( .A(n464), .Z(n388) );
  GTECH_NAND3 U438 ( .A(n10), .B(n465), .C(N155), .Z(n464) );
  GTECH_NAND2 U439 ( .A(n466), .B(N155), .Z(n456) );
  GTECH_XOR2 U440 ( .A(n463), .B(n28), .Z(n466) );
  GTECH_AND2 U441 ( .A(N155), .B(n467), .Z(N134) );
  GTECH_NOT U442 ( .A(n13), .Z(n467) );
  GTECH_AND2 U443 ( .A(N155), .B(n468), .Z(N133) );
  GTECH_NOT U444 ( .A(n14), .Z(n468) );
  GTECH_AND2 U445 ( .A(N155), .B(n469), .Z(N132) );
  GTECH_NOT U446 ( .A(n15), .Z(n469) );
  GTECH_AND2 U447 ( .A(N155), .B(n470), .Z(N131) );
  GTECH_NOT U448 ( .A(n16), .Z(n470) );
  GTECH_AND2 U449 ( .A(N155), .B(n471), .Z(N130) );
  GTECH_NOT U450 ( .A(n17), .Z(n471) );
  GTECH_AND2 U451 ( .A(N155), .B(n472), .Z(N129) );
  GTECH_NOT U452 ( .A(n18), .Z(n472) );
  GTECH_AND2 U453 ( .A(N155), .B(n473), .Z(N128) );
  GTECH_NOT U454 ( .A(n19), .Z(n473) );
  GTECH_AND2 U455 ( .A(N155), .B(n474), .Z(N127) );
  GTECH_NOT U456 ( .A(n20), .Z(n474) );
  GTECH_AND2 U457 ( .A(N155), .B(n475), .Z(N126) );
  GTECH_NOT U458 ( .A(n21), .Z(n475) );
  GTECH_AND2 U459 ( .A(N155), .B(n476), .Z(N125) );
  GTECH_NOT U460 ( .A(n22), .Z(n476) );
  GTECH_AND2 U461 ( .A(N155), .B(n477), .Z(N124) );
  GTECH_NOT U462 ( .A(n23), .Z(n477) );
  GTECH_AND2 U463 ( .A(N155), .B(n478), .Z(N123) );
  GTECH_NOT U464 ( .A(n24), .Z(n478) );
  GTECH_AND2 U465 ( .A(N155), .B(n479), .Z(N122) );
  GTECH_NOT U466 ( .A(n25), .Z(n479) );
  GTECH_AND2 U467 ( .A(N155), .B(n480), .Z(N121) );
  GTECH_NOT U468 ( .A(n26), .Z(n480) );
  GTECH_AND2 U469 ( .A(N155), .B(n481), .Z(N120) );
  GTECH_NOT U470 ( .A(n27), .Z(n481) );
  GTECH_NOT U471 ( .A(n390), .Z(N155) );
  GTECH_NAND4 U472 ( .A(n8), .B(n7), .C(n9), .D(n482), .Z(n390) );
  GTECH_AND3 U473 ( .A(n377), .B(n398), .C(n6), .Z(n482) );
  GTECH_NOT U474 ( .A(n338), .Z(n398) );
  GTECH_NOT U475 ( .A(n483), .Z(N116) );
  GTECH_AOI222 U476 ( .A(n359), .B(n387), .C(n361), .D(n389), .E(n385), .F(
        n357), .Z(n483) );
  GTECH_XOR2 U477 ( .A(n484), .B(n485), .Z(n385) );
  GTECH_ADD_ABC U478 ( .A(n354), .B(n31), .C(n486), .COUT(n485) );
  GTECH_XOR2 U479 ( .A(n487), .B(n484), .Z(n389) );
  GTECH_XOR2 U480 ( .A(n387), .B(n355), .Z(n484) );
  GTECH_NAND2 U481 ( .A(n488), .B(n489), .Z(n487) );
  GTECH_OAI21 U482 ( .A(n354), .B(n393), .C(n490), .Z(n489) );
  GTECH_OR_NOT U483 ( .A(n31), .B(n354), .Z(n488) );
  GTECH_NOT U484 ( .A(n30), .Z(n387) );
  GTECH_NAND2 U485 ( .A(n370), .B(n491), .Z(N115) );
  GTECH_NOT U486 ( .A(N41), .Z(n491) );
  GTECH_NAND2 U487 ( .A(n377), .B(n371), .Z(N41) );
  GTECH_NAND2 U488 ( .A(Ld), .B(n377), .Z(n371) );
  GTECH_NOT U489 ( .A(n492), .Z(N113) );
  GTECH_AOI222 U490 ( .A(n359), .B(n393), .C(n361), .D(n394), .E(n392), .F(
        n357), .Z(n492) );
  GTECH_XOR2 U491 ( .A(n493), .B(n486), .Z(n392) );
  GTECH_ADD_ABC U492 ( .A(n353), .B(n32), .C(n494), .COUT(n486) );
  GTECH_NOT U493 ( .A(n495), .Z(n394) );
  GTECH_XOR2 U494 ( .A(n493), .B(n496), .Z(n495) );
  GTECH_NOT U495 ( .A(n490), .Z(n496) );
  GTECH_OAI21 U496 ( .A(n32), .B(n497), .C(n498), .Z(n490) );
  GTECH_OAI21 U497 ( .A(n353), .B(n401), .C(n499), .Z(n498) );
  GTECH_NOT U498 ( .A(n353), .Z(n497) );
  GTECH_XOR2 U499 ( .A(n393), .B(n354), .Z(n493) );
  GTECH_NOT U500 ( .A(n31), .Z(n393) );
  GTECH_NOT U501 ( .A(n500), .Z(N112) );
  GTECH_AOI222 U502 ( .A(n359), .B(n401), .C(n361), .D(n402), .E(n400), .F(
        n357), .Z(n500) );
  GTECH_XOR2 U503 ( .A(n501), .B(n494), .Z(n400) );
  GTECH_ADD_ABC U504 ( .A(n33), .B(n352), .C(n502), .COUT(n494) );
  GTECH_NOT U505 ( .A(n503), .Z(n402) );
  GTECH_XOR2 U506 ( .A(n501), .B(n504), .Z(n503) );
  GTECH_NOT U507 ( .A(n499), .Z(n504) );
  GTECH_OAI21 U508 ( .A(n33), .B(n505), .C(n506), .Z(n499) );
  GTECH_OAI21 U509 ( .A(n352), .B(n405), .C(n507), .Z(n506) );
  GTECH_XOR2 U510 ( .A(n401), .B(n353), .Z(n501) );
  GTECH_NOT U511 ( .A(n32), .Z(n401) );
  GTECH_NOT U512 ( .A(n508), .Z(N111) );
  GTECH_AOI222 U513 ( .A(n359), .B(n405), .C(n361), .D(n406), .E(n404), .F(
        n357), .Z(n508) );
  GTECH_XOR2 U514 ( .A(n509), .B(n502), .Z(n404) );
  GTECH_ADD_ABC U515 ( .A(n34), .B(n351), .C(n510), .COUT(n502) );
  GTECH_NOT U516 ( .A(n511), .Z(n406) );
  GTECH_XOR2 U517 ( .A(n509), .B(n512), .Z(n511) );
  GTECH_NOT U518 ( .A(n507), .Z(n512) );
  GTECH_OAI21 U519 ( .A(n34), .B(n513), .C(n514), .Z(n507) );
  GTECH_OAI21 U520 ( .A(n351), .B(n409), .C(n515), .Z(n514) );
  GTECH_XOR2 U521 ( .A(n505), .B(n33), .Z(n509) );
  GTECH_NOT U522 ( .A(n352), .Z(n505) );
  GTECH_NOT U523 ( .A(n33), .Z(n405) );
  GTECH_NOT U524 ( .A(n516), .Z(N110) );
  GTECH_AOI222 U525 ( .A(n359), .B(n409), .C(n361), .D(n410), .E(n408), .F(
        n357), .Z(n516) );
  GTECH_XOR2 U526 ( .A(n517), .B(n510), .Z(n408) );
  GTECH_ADD_ABC U527 ( .A(n35), .B(n350), .C(n518), .COUT(n510) );
  GTECH_NOT U528 ( .A(n519), .Z(n410) );
  GTECH_XOR2 U529 ( .A(n517), .B(n520), .Z(n519) );
  GTECH_NOT U530 ( .A(n515), .Z(n520) );
  GTECH_OAI21 U531 ( .A(n35), .B(n521), .C(n522), .Z(n515) );
  GTECH_OAI21 U532 ( .A(n350), .B(n413), .C(n523), .Z(n522) );
  GTECH_XOR2 U533 ( .A(n513), .B(n34), .Z(n517) );
  GTECH_NOT U534 ( .A(n351), .Z(n513) );
  GTECH_NOT U535 ( .A(n34), .Z(n409) );
  GTECH_NOT U536 ( .A(n524), .Z(N109) );
  GTECH_AOI222 U537 ( .A(n359), .B(n413), .C(n361), .D(n414), .E(n412), .F(
        n357), .Z(n524) );
  GTECH_XOR2 U538 ( .A(n525), .B(n518), .Z(n412) );
  GTECH_ADD_ABC U539 ( .A(n36), .B(n349), .C(n526), .COUT(n518) );
  GTECH_NOT U540 ( .A(n527), .Z(n414) );
  GTECH_XOR2 U541 ( .A(n525), .B(n528), .Z(n527) );
  GTECH_NOT U542 ( .A(n523), .Z(n528) );
  GTECH_OAI21 U543 ( .A(n36), .B(n529), .C(n530), .Z(n523) );
  GTECH_OAI21 U544 ( .A(n349), .B(n417), .C(n531), .Z(n530) );
  GTECH_XOR2 U545 ( .A(n521), .B(n35), .Z(n525) );
  GTECH_NOT U546 ( .A(n350), .Z(n521) );
  GTECH_NOT U547 ( .A(n35), .Z(n413) );
  GTECH_NOT U548 ( .A(n532), .Z(N108) );
  GTECH_AOI222 U549 ( .A(n359), .B(n417), .C(n361), .D(n418), .E(n416), .F(
        n357), .Z(n532) );
  GTECH_XOR2 U550 ( .A(n533), .B(n526), .Z(n416) );
  GTECH_ADD_ABC U551 ( .A(n37), .B(n348), .C(n534), .COUT(n526) );
  GTECH_NOT U552 ( .A(n535), .Z(n418) );
  GTECH_XOR2 U553 ( .A(n533), .B(n536), .Z(n535) );
  GTECH_NOT U554 ( .A(n531), .Z(n536) );
  GTECH_OAI21 U555 ( .A(n37), .B(n537), .C(n538), .Z(n531) );
  GTECH_OAI21 U556 ( .A(n348), .B(n421), .C(n539), .Z(n538) );
  GTECH_XOR2 U557 ( .A(n529), .B(n36), .Z(n533) );
  GTECH_NOT U558 ( .A(n349), .Z(n529) );
  GTECH_NOT U559 ( .A(n36), .Z(n417) );
  GTECH_NOT U560 ( .A(n540), .Z(N107) );
  GTECH_AOI222 U561 ( .A(n359), .B(n421), .C(n361), .D(n422), .E(n420), .F(
        n357), .Z(n540) );
  GTECH_XOR2 U562 ( .A(n541), .B(n534), .Z(n420) );
  GTECH_ADD_ABC U563 ( .A(n38), .B(n347), .C(n542), .COUT(n534) );
  GTECH_NOT U564 ( .A(n543), .Z(n422) );
  GTECH_XOR2 U565 ( .A(n541), .B(n544), .Z(n543) );
  GTECH_NOT U566 ( .A(n539), .Z(n544) );
  GTECH_OAI21 U567 ( .A(n38), .B(n545), .C(n546), .Z(n539) );
  GTECH_OAI21 U568 ( .A(n347), .B(n425), .C(n547), .Z(n546) );
  GTECH_XOR2 U569 ( .A(n537), .B(n37), .Z(n541) );
  GTECH_NOT U570 ( .A(n348), .Z(n537) );
  GTECH_NOT U571 ( .A(n37), .Z(n421) );
  GTECH_NOT U572 ( .A(n548), .Z(N106) );
  GTECH_AOI222 U573 ( .A(n359), .B(n425), .C(n361), .D(n426), .E(n424), .F(
        n357), .Z(n548) );
  GTECH_XOR2 U574 ( .A(n549), .B(n542), .Z(n424) );
  GTECH_ADD_ABC U575 ( .A(n39), .B(n346), .C(n550), .COUT(n542) );
  GTECH_NOT U576 ( .A(n551), .Z(n426) );
  GTECH_XOR2 U577 ( .A(n549), .B(n552), .Z(n551) );
  GTECH_NOT U578 ( .A(n547), .Z(n552) );
  GTECH_OAI21 U579 ( .A(n39), .B(n553), .C(n554), .Z(n547) );
  GTECH_OAI21 U580 ( .A(n346), .B(n429), .C(n555), .Z(n554) );
  GTECH_XOR2 U581 ( .A(n545), .B(n38), .Z(n549) );
  GTECH_NOT U582 ( .A(n347), .Z(n545) );
  GTECH_NOT U583 ( .A(n38), .Z(n425) );
  GTECH_NOT U584 ( .A(n556), .Z(N105) );
  GTECH_AOI222 U585 ( .A(n359), .B(n429), .C(n361), .D(n430), .E(n428), .F(
        n357), .Z(n556) );
  GTECH_XOR2 U586 ( .A(n557), .B(n550), .Z(n428) );
  GTECH_ADD_ABC U587 ( .A(n40), .B(n345), .C(n558), .COUT(n550) );
  GTECH_NOT U588 ( .A(n559), .Z(n430) );
  GTECH_XOR2 U589 ( .A(n557), .B(n560), .Z(n559) );
  GTECH_NOT U590 ( .A(n555), .Z(n560) );
  GTECH_OAI21 U591 ( .A(n40), .B(n561), .C(n562), .Z(n555) );
  GTECH_OAI21 U592 ( .A(n345), .B(n433), .C(n563), .Z(n562) );
  GTECH_XOR2 U593 ( .A(n553), .B(n39), .Z(n557) );
  GTECH_NOT U594 ( .A(n346), .Z(n553) );
  GTECH_NOT U595 ( .A(n39), .Z(n429) );
  GTECH_NOT U596 ( .A(n564), .Z(N104) );
  GTECH_AOI222 U597 ( .A(n359), .B(n433), .C(n361), .D(n434), .E(n432), .F(
        n357), .Z(n564) );
  GTECH_XOR2 U598 ( .A(n565), .B(n558), .Z(n432) );
  GTECH_ADD_ABC U599 ( .A(n41), .B(n344), .C(n566), .COUT(n558) );
  GTECH_NOT U600 ( .A(n567), .Z(n434) );
  GTECH_XOR2 U601 ( .A(n565), .B(n568), .Z(n567) );
  GTECH_NOT U602 ( .A(n563), .Z(n568) );
  GTECH_OAI21 U603 ( .A(n41), .B(n569), .C(n570), .Z(n563) );
  GTECH_OAI21 U604 ( .A(n344), .B(n437), .C(n571), .Z(n570) );
  GTECH_XOR2 U605 ( .A(n561), .B(n40), .Z(n565) );
  GTECH_NOT U606 ( .A(n345), .Z(n561) );
  GTECH_NOT U607 ( .A(n40), .Z(n433) );
  GTECH_NOT U608 ( .A(n572), .Z(N103) );
  GTECH_AOI222 U609 ( .A(n359), .B(n437), .C(n361), .D(n438), .E(n436), .F(
        n357), .Z(n572) );
  GTECH_XOR2 U610 ( .A(n573), .B(n566), .Z(n436) );
  GTECH_ADD_ABC U611 ( .A(n42), .B(n343), .C(n574), .COUT(n566) );
  GTECH_NOT U612 ( .A(n575), .Z(n438) );
  GTECH_XOR2 U613 ( .A(n573), .B(n576), .Z(n575) );
  GTECH_NOT U614 ( .A(n571), .Z(n576) );
  GTECH_OAI21 U615 ( .A(n42), .B(n577), .C(n578), .Z(n571) );
  GTECH_OAI21 U616 ( .A(n343), .B(n441), .C(n579), .Z(n578) );
  GTECH_XOR2 U617 ( .A(n569), .B(n41), .Z(n573) );
  GTECH_NOT U618 ( .A(n344), .Z(n569) );
  GTECH_NOT U619 ( .A(n41), .Z(n437) );
  GTECH_NOT U620 ( .A(n580), .Z(N102) );
  GTECH_AOI222 U621 ( .A(n359), .B(n441), .C(n361), .D(n442), .E(n440), .F(
        n357), .Z(n580) );
  GTECH_XOR2 U622 ( .A(n581), .B(n574), .Z(n440) );
  GTECH_ADD_ABC U623 ( .A(n43), .B(n342), .C(n582), .COUT(n574) );
  GTECH_NOT U624 ( .A(n583), .Z(n442) );
  GTECH_XOR2 U625 ( .A(n581), .B(n584), .Z(n583) );
  GTECH_NOT U626 ( .A(n579), .Z(n584) );
  GTECH_OAI21 U627 ( .A(n43), .B(n585), .C(n586), .Z(n579) );
  GTECH_OAI21 U628 ( .A(n342), .B(n445), .C(n587), .Z(n586) );
  GTECH_XOR2 U629 ( .A(n577), .B(n42), .Z(n581) );
  GTECH_NOT U630 ( .A(n343), .Z(n577) );
  GTECH_NOT U631 ( .A(n42), .Z(n441) );
  GTECH_NOT U632 ( .A(n588), .Z(N101) );
  GTECH_AOI222 U633 ( .A(n359), .B(n445), .C(n361), .D(n446), .E(n444), .F(
        n357), .Z(n588) );
  GTECH_XOR2 U634 ( .A(n589), .B(n582), .Z(n444) );
  GTECH_ADD_ABC U635 ( .A(n29), .B(n341), .C(n590), .COUT(n582) );
  GTECH_NOT U636 ( .A(n591), .Z(n446) );
  GTECH_XOR2 U637 ( .A(n589), .B(n592), .Z(n591) );
  GTECH_NOT U638 ( .A(n587), .Z(n592) );
  GTECH_OAI21 U639 ( .A(n29), .B(n593), .C(n594), .Z(n587) );
  GTECH_OAI21 U640 ( .A(n341), .B(n449), .C(n595), .Z(n594) );
  GTECH_XOR2 U641 ( .A(n585), .B(n43), .Z(n589) );
  GTECH_NOT U642 ( .A(n342), .Z(n585) );
  GTECH_NOT U643 ( .A(n43), .Z(n445) );
  GTECH_NOT U644 ( .A(n596), .Z(N100) );
  GTECH_AOI222 U645 ( .A(n448), .B(n357), .C(n359), .D(n449), .E(n361), .F(
        n450), .Z(n596) );
  GTECH_NOT U646 ( .A(n597), .Z(n450) );
  GTECH_XOR2 U647 ( .A(n598), .B(n599), .Z(n597) );
  GTECH_NOT U648 ( .A(n595), .Z(n599) );
  GTECH_OAI21 U649 ( .A(n11), .B(n600), .C(n601), .Z(n595) );
  GTECH_OAI21 U650 ( .A(n340), .B(n360), .C(n455), .Z(n601) );
  GTECH_NAND2 U651 ( .A(n12), .B(n461), .Z(n455) );
  GTECH_NOT U652 ( .A(n11), .Z(n360) );
  GTECH_NOT U653 ( .A(n340), .Z(n600) );
  GTECH_NOT U654 ( .A(n369), .Z(n361) );
  GTECH_NAND2 U655 ( .A(N82), .B(n10), .Z(n369) );
  GTECH_NOT U656 ( .A(n602), .Z(N82) );
  GTECH_NOT U657 ( .A(n29), .Z(n449) );
  GTECH_OAI21 U658 ( .A(n10), .B(n602), .C(n603), .Z(n359) );
  GTECH_NAND3 U659 ( .A(n28), .B(n375), .C(n10), .Z(n603) );
  GTECH_NAND2 U660 ( .A(n375), .B(n465), .Z(n602) );
  GTECH_NOT U661 ( .A(n28), .Z(n465) );
  GTECH_NOT U662 ( .A(n368), .Z(n357) );
  GTECH_NAND3 U663 ( .A(n375), .B(n463), .C(n28), .Z(n368) );
  GTECH_NOT U664 ( .A(n10), .Z(n463) );
  GTECH_NOT U665 ( .A(n370), .Z(n375) );
  GTECH_OAI21 U666 ( .A(n373), .B(n374), .C(n604), .Z(n370) );
  GTECH_AND2 U667 ( .A(n376), .B(n377), .Z(n604) );
  GTECH_NOT U668 ( .A(Rst), .Z(n377) );
  GTECH_NOT U669 ( .A(Ld), .Z(n376) );
  GTECH_NOT U670 ( .A(n9), .Z(n374) );
  GTECH_NAND2 U671 ( .A(n8), .B(n379), .Z(n373) );
  GTECH_NOT U672 ( .A(n382), .Z(n379) );
  GTECH_NAND2 U673 ( .A(n7), .B(n381), .Z(n382) );
  GTECH_NOT U674 ( .A(n605), .Z(n381) );
  GTECH_NAND2 U675 ( .A(n6), .B(n338), .Z(n605) );
  GTECH_XOR2 U676 ( .A(n598), .B(n590), .Z(n448) );
  GTECH_ADD_ABC U677 ( .A(n340), .B(n11), .C(n459), .COUT(n590) );
  GTECH_NAND2 U678 ( .A(n364), .B(n461), .Z(n459) );
  GTECH_NOT U679 ( .A(n339), .Z(n461) );
  GTECH_NOT U680 ( .A(n12), .Z(n364) );
  GTECH_XOR2 U681 ( .A(n593), .B(n29), .Z(n598) );
  GTECH_NOT U682 ( .A(n341), .Z(n593) );
endmodule

