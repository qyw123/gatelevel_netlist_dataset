
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138;

  GTECH_XOR2 U91 ( .A(n72), .B(n73), .Z(sum[9]) );
  GTECH_XNOR2 U92 ( .A(n74), .B(n75), .Z(sum[8]) );
  GTECH_XNOR2 U93 ( .A(n76), .B(n77), .Z(sum[7]) );
  GTECH_AOI21 U94 ( .A(n78), .B(n79), .C(n80), .Z(n77) );
  GTECH_XOR2 U95 ( .A(n79), .B(n78), .Z(sum[6]) );
  GTECH_AO22 U96 ( .A(b[5]), .B(a[5]), .C(n81), .D(n82), .Z(n78) );
  GTECH_XOR2 U97 ( .A(n82), .B(n81), .Z(sum[5]) );
  GTECH_AO21 U98 ( .A(n83), .B(n84), .C(n85), .Z(n81) );
  GTECH_XOR2 U99 ( .A(n84), .B(n83), .Z(sum[4]) );
  GTECH_XNOR2 U100 ( .A(n86), .B(n87), .Z(sum[3]) );
  GTECH_AOI21 U101 ( .A(n88), .B(n89), .C(n90), .Z(n87) );
  GTECH_XOR2 U102 ( .A(n89), .B(n88), .Z(sum[2]) );
  GTECH_AO22 U103 ( .A(b[1]), .B(a[1]), .C(n91), .D(n92), .Z(n88) );
  GTECH_XOR2 U104 ( .A(n92), .B(n91), .Z(sum[1]) );
  GTECH_AO22 U105 ( .A(n93), .B(cin), .C(a[0]), .D(b[0]), .Z(n91) );
  GTECH_XNOR2 U106 ( .A(n94), .B(n95), .Z(sum[15]) );
  GTECH_AOI21 U107 ( .A(n96), .B(n97), .C(n98), .Z(n95) );
  GTECH_XOR2 U108 ( .A(n97), .B(n96), .Z(sum[14]) );
  GTECH_AO22 U109 ( .A(b[13]), .B(a[13]), .C(n99), .D(n100), .Z(n96) );
  GTECH_XOR2 U110 ( .A(n100), .B(n99), .Z(sum[13]) );
  GTECH_AO21 U111 ( .A(cout), .B(n101), .C(n102), .Z(n99) );
  GTECH_XOR2 U112 ( .A(cout), .B(n101), .Z(sum[12]) );
  GTECH_XNOR2 U113 ( .A(n103), .B(n104), .Z(sum[11]) );
  GTECH_AOI21 U114 ( .A(n105), .B(n106), .C(n107), .Z(n104) );
  GTECH_XOR2 U115 ( .A(n106), .B(n105), .Z(sum[10]) );
  GTECH_AO22 U116 ( .A(b[9]), .B(a[9]), .C(n73), .D(n72), .Z(n105) );
  GTECH_AO22 U117 ( .A(a[8]), .B(b[8]), .C(n108), .D(n74), .Z(n73) );
  GTECH_NOT U118 ( .A(n75), .Z(n108) );
  GTECH_XNOR2 U119 ( .A(n109), .B(n93), .Z(sum[0]) );
  GTECH_OAI21 U120 ( .A(n75), .B(n110), .C(n111), .Z(cout) );
  GTECH_OA21 U121 ( .A(n112), .B(n113), .C(n114), .Z(n75) );
  GTECH_NOT U122 ( .A(n83), .Z(n112) );
  GTECH_OAI21 U123 ( .A(n115), .B(n109), .C(n116), .Z(n83) );
  GTECH_NOT U124 ( .A(cin), .Z(n109) );
  GTECH_NOR3 U125 ( .A(n113), .B(n115), .C(n110), .Z(Pm) );
  GTECH_NAND5 U126 ( .A(n89), .B(n92), .C(n86), .D(n117), .E(n93), .Z(n115) );
  GTECH_XOR2 U127 ( .A(a[0]), .B(b[0]), .Z(n93) );
  GTECH_OAI21 U128 ( .A(n118), .B(n110), .C(n111), .Z(Gm) );
  GTECH_AOI2N2 U129 ( .A(b[15]), .B(a[15]), .C(n119), .D(n120), .Z(n111) );
  GTECH_NOT U130 ( .A(n94), .Z(n120) );
  GTECH_AOI21 U131 ( .A(n121), .B(n97), .C(n98), .Z(n119) );
  GTECH_AND2 U132 ( .A(b[14]), .B(a[14]), .Z(n98) );
  GTECH_AO22 U133 ( .A(n100), .B(n102), .C(b[13]), .D(a[13]), .Z(n121) );
  GTECH_NAND4 U134 ( .A(n101), .B(n94), .C(n97), .D(n100), .Z(n110) );
  GTECH_XOR2 U135 ( .A(a[13]), .B(b[13]), .Z(n100) );
  GTECH_XOR2 U136 ( .A(a[14]), .B(b[14]), .Z(n97) );
  GTECH_XOR2 U137 ( .A(a[15]), .B(b[15]), .Z(n94) );
  GTECH_OA21 U138 ( .A(b[12]), .B(a[12]), .C(n122), .Z(n101) );
  GTECH_NOT U139 ( .A(n102), .Z(n122) );
  GTECH_AND2 U140 ( .A(b[12]), .B(a[12]), .Z(n102) );
  GTECH_OA21 U141 ( .A(n116), .B(n113), .C(n114), .Z(n118) );
  GTECH_AOI2N2 U142 ( .A(b[11]), .B(a[11]), .C(n123), .D(n124), .Z(n114) );
  GTECH_NOT U143 ( .A(n103), .Z(n124) );
  GTECH_AOI21 U144 ( .A(n125), .B(n106), .C(n107), .Z(n123) );
  GTECH_AND2 U145 ( .A(a[10]), .B(b[10]), .Z(n107) );
  GTECH_OAI21 U146 ( .A(n126), .B(n127), .C(n128), .Z(n125) );
  GTECH_NAND3 U147 ( .A(a[8]), .B(n72), .C(b[8]), .Z(n128) );
  GTECH_NAND4 U148 ( .A(n74), .B(n103), .C(n106), .D(n72), .Z(n113) );
  GTECH_XOR2 U149 ( .A(n127), .B(n126), .Z(n72) );
  GTECH_NOT U150 ( .A(b[9]), .Z(n126) );
  GTECH_NOT U151 ( .A(a[9]), .Z(n127) );
  GTECH_XOR2 U152 ( .A(a[10]), .B(b[10]), .Z(n106) );
  GTECH_XOR2 U153 ( .A(a[11]), .B(b[11]), .Z(n103) );
  GTECH_XOR2 U154 ( .A(a[8]), .B(b[8]), .Z(n74) );
  GTECH_AOI222 U155 ( .A(n117), .B(n129), .C(b[7]), .D(a[7]), .E(n76), .F(n130), .Z(n116) );
  GTECH_AO21 U156 ( .A(n131), .B(n79), .C(n80), .Z(n130) );
  GTECH_AND2 U157 ( .A(b[6]), .B(a[6]), .Z(n80) );
  GTECH_AO22 U158 ( .A(n82), .B(n85), .C(b[5]), .D(a[5]), .Z(n131) );
  GTECH_OAI2N2 U159 ( .A(n132), .B(n133), .C(b[3]), .D(a[3]), .Z(n129) );
  GTECH_NOT U160 ( .A(n86), .Z(n133) );
  GTECH_XOR2 U161 ( .A(a[3]), .B(b[3]), .Z(n86) );
  GTECH_AOI21 U162 ( .A(n134), .B(n89), .C(n90), .Z(n132) );
  GTECH_AND2 U163 ( .A(b[2]), .B(a[2]), .Z(n90) );
  GTECH_XOR2 U164 ( .A(a[2]), .B(b[2]), .Z(n89) );
  GTECH_OAI21 U165 ( .A(n135), .B(n136), .C(n137), .Z(n134) );
  GTECH_NAND3 U166 ( .A(a[0]), .B(n92), .C(b[0]), .Z(n137) );
  GTECH_XOR2 U167 ( .A(n136), .B(n135), .Z(n92) );
  GTECH_NOT U168 ( .A(a[1]), .Z(n136) );
  GTECH_NOT U169 ( .A(b[1]), .Z(n135) );
  GTECH_AND4 U170 ( .A(n84), .B(n82), .C(n79), .D(n76), .Z(n117) );
  GTECH_XOR2 U171 ( .A(a[7]), .B(b[7]), .Z(n76) );
  GTECH_XOR2 U172 ( .A(a[6]), .B(b[6]), .Z(n79) );
  GTECH_XOR2 U173 ( .A(a[5]), .B(b[5]), .Z(n82) );
  GTECH_OA21 U174 ( .A(b[4]), .B(a[4]), .C(n138), .Z(n84) );
  GTECH_NOT U175 ( .A(n85), .Z(n138) );
  GTECH_AND2 U176 ( .A(b[4]), .B(a[4]), .Z(n85) );
endmodule

