
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_OR_NOT U83 ( .A(n97), .B(n93), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n98), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n98) );
  GTECH_OAI21 U86 ( .A(n99), .B(n100), .C(n101), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  GTECH_NOT U88 ( .A(n103), .Z(n99) );
  GTECH_OR_NOT U89 ( .A(n105), .B(I_b[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n106), .Z(n84) );
  GTECH_OR_NOT U91 ( .A(n107), .B(n108), .Z(n106) );
  GTECH_XOR2 U92 ( .A(n109), .B(n108), .Z(N153) );
  GTECH_NOT U93 ( .A(n110), .Z(n108) );
  GTECH_XOR3 U94 ( .A(n97), .B(n93), .C(n95), .Z(n110) );
  GTECH_XOR3 U95 ( .A(n102), .B(n104), .C(n103), .Z(n95) );
  GTECH_OAI21 U96 ( .A(n111), .B(n112), .C(n113), .Z(n103) );
  GTECH_OAI21 U97 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_NOT U98 ( .A(n115), .Z(n111) );
  GTECH_NOT U99 ( .A(n117), .Z(n104) );
  GTECH_OR_NOT U100 ( .A(n118), .B(I_b[7]), .Z(n117) );
  GTECH_NOT U101 ( .A(n100), .Z(n102) );
  GTECH_OR_NOT U102 ( .A(n119), .B(I_a[7]), .Z(n100) );
  GTECH_NOT U103 ( .A(I_b[6]), .Z(n119) );
  GTECH_ADD_ABC U104 ( .A(n120), .B(n121), .C(n122), .COUT(n93) );
  GTECH_NOT U105 ( .A(n123), .Z(n122) );
  GTECH_XOR2 U106 ( .A(n124), .B(n125), .Z(n121) );
  GTECH_AND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n125) );
  GTECH_NOT U108 ( .A(n94), .Z(n97) );
  GTECH_OR_NOT U109 ( .A(n124), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U110 ( .A(n107), .Z(n109) );
  GTECH_OR_NOT U111 ( .A(n126), .B(n127), .Z(n107) );
  GTECH_XOR2 U112 ( .A(n126), .B(n128), .Z(N152) );
  GTECH_NOT U113 ( .A(n127), .Z(n128) );
  GTECH_XOR4 U114 ( .A(n129), .B(n124), .C(n120), .D(n123), .Z(n127) );
  GTECH_XOR3 U115 ( .A(n114), .B(n116), .C(n115), .Z(n123) );
  GTECH_OAI21 U116 ( .A(n130), .B(n131), .C(n132), .Z(n115) );
  GTECH_OAI21 U117 ( .A(n133), .B(n134), .C(n135), .Z(n132) );
  GTECH_NOT U118 ( .A(n134), .Z(n130) );
  GTECH_NOT U119 ( .A(n136), .Z(n116) );
  GTECH_OR_NOT U120 ( .A(n137), .B(I_b[7]), .Z(n136) );
  GTECH_NOT U121 ( .A(n112), .Z(n114) );
  GTECH_OR_NOT U122 ( .A(n118), .B(I_b[6]), .Z(n112) );
  GTECH_NOT U123 ( .A(I_a[6]), .Z(n118) );
  GTECH_ADD_ABC U124 ( .A(n138), .B(n139), .C(n140), .COUT(n120) );
  GTECH_NOT U125 ( .A(n141), .Z(n140) );
  GTECH_XOR3 U126 ( .A(n142), .B(n143), .C(n144), .Z(n139) );
  GTECH_OA21 U127 ( .A(n144), .B(n145), .C(n146), .Z(n124) );
  GTECH_OAI21 U128 ( .A(n142), .B(n147), .C(n143), .Z(n146) );
  GTECH_NOT U129 ( .A(n145), .Z(n142) );
  GTECH_NOT U130 ( .A(n147), .Z(n144) );
  GTECH_AND2 U131 ( .A(I_b[5]), .B(I_a[7]), .Z(n129) );
  GTECH_ADD_ABC U132 ( .A(n148), .B(n149), .C(n150), .COUT(n126) );
  GTECH_NOT U133 ( .A(n151), .Z(n150) );
  GTECH_OA22 U134 ( .A(n152), .B(n105), .C(n153), .D(n154), .Z(n149) );
  GTECH_OA21 U135 ( .A(n155), .B(n156), .C(n157), .Z(n148) );
  GTECH_XOR3 U136 ( .A(n158), .B(n151), .C(n159), .Z(N151) );
  GTECH_OA21 U137 ( .A(n155), .B(n156), .C(n157), .Z(n159) );
  GTECH_OAI21 U138 ( .A(n160), .B(n161), .C(n162), .Z(n157) );
  GTECH_XOR2 U139 ( .A(n163), .B(n138), .Z(n151) );
  GTECH_ADD_ABC U140 ( .A(n164), .B(n165), .C(n166), .COUT(n138) );
  GTECH_NOT U141 ( .A(n167), .Z(n166) );
  GTECH_XOR3 U142 ( .A(n168), .B(n169), .C(n170), .Z(n165) );
  GTECH_XOR4 U143 ( .A(n143), .B(n147), .C(n145), .D(n141), .Z(n163) );
  GTECH_XOR3 U144 ( .A(n133), .B(n135), .C(n134), .Z(n141) );
  GTECH_OAI21 U145 ( .A(n171), .B(n172), .C(n173), .Z(n134) );
  GTECH_OAI21 U146 ( .A(n174), .B(n175), .C(n176), .Z(n173) );
  GTECH_NOT U147 ( .A(n175), .Z(n171) );
  GTECH_NOT U148 ( .A(n177), .Z(n135) );
  GTECH_OR_NOT U149 ( .A(n178), .B(I_b[7]), .Z(n177) );
  GTECH_NOT U150 ( .A(n131), .Z(n133) );
  GTECH_OR_NOT U151 ( .A(n137), .B(I_b[6]), .Z(n131) );
  GTECH_NOT U152 ( .A(I_a[5]), .Z(n137) );
  GTECH_OR_NOT U153 ( .A(n179), .B(I_a[7]), .Z(n145) );
  GTECH_OAI21 U154 ( .A(n170), .B(n180), .C(n181), .Z(n147) );
  GTECH_OAI21 U155 ( .A(n168), .B(n182), .C(n169), .Z(n181) );
  GTECH_NOT U156 ( .A(n180), .Z(n168) );
  GTECH_NOT U157 ( .A(n182), .Z(n170) );
  GTECH_NOT U158 ( .A(n183), .Z(n143) );
  GTECH_OR_NOT U159 ( .A(n184), .B(I_a[6]), .Z(n183) );
  GTECH_OA22 U160 ( .A(n152), .B(n105), .C(n153), .D(n154), .Z(n158) );
  GTECH_NOT U161 ( .A(n185), .Z(n154) );
  GTECH_NOT U162 ( .A(I_a[7]), .Z(n105) );
  GTECH_XOR3 U163 ( .A(n155), .B(n160), .C(n186), .Z(N150) );
  GTECH_NOT U164 ( .A(n162), .Z(n186) );
  GTECH_XOR2 U165 ( .A(n187), .B(n164), .Z(n162) );
  GTECH_ADD_ABC U166 ( .A(n188), .B(n189), .C(n190), .COUT(n164) );
  GTECH_NOT U167 ( .A(n191), .Z(n190) );
  GTECH_XOR3 U168 ( .A(n192), .B(n193), .C(n194), .Z(n189) );
  GTECH_XOR4 U169 ( .A(n169), .B(n182), .C(n180), .D(n167), .Z(n187) );
  GTECH_XOR3 U170 ( .A(n174), .B(n176), .C(n175), .Z(n167) );
  GTECH_OAI21 U171 ( .A(n195), .B(n196), .C(n197), .Z(n175) );
  GTECH_OAI21 U172 ( .A(n198), .B(n199), .C(n200), .Z(n197) );
  GTECH_NOT U173 ( .A(n199), .Z(n195) );
  GTECH_NOT U174 ( .A(n201), .Z(n176) );
  GTECH_OR_NOT U175 ( .A(n202), .B(I_b[7]), .Z(n201) );
  GTECH_NOT U176 ( .A(n172), .Z(n174) );
  GTECH_OR_NOT U177 ( .A(n178), .B(I_b[6]), .Z(n172) );
  GTECH_OR_NOT U178 ( .A(n179), .B(I_a[6]), .Z(n180) );
  GTECH_OAI21 U179 ( .A(n194), .B(n203), .C(n204), .Z(n182) );
  GTECH_OAI21 U180 ( .A(n192), .B(n205), .C(n193), .Z(n204) );
  GTECH_NOT U181 ( .A(n203), .Z(n192) );
  GTECH_NOT U182 ( .A(n205), .Z(n194) );
  GTECH_NOT U183 ( .A(n206), .Z(n169) );
  GTECH_OR_NOT U184 ( .A(n184), .B(I_a[5]), .Z(n206) );
  GTECH_NOT U185 ( .A(I_b[5]), .Z(n184) );
  GTECH_NOT U186 ( .A(n156), .Z(n160) );
  GTECH_XOR2 U187 ( .A(n185), .B(n153), .Z(n156) );
  GTECH_NOT U188 ( .A(n207), .Z(n153) );
  GTECH_OAI2N2 U189 ( .A(n208), .B(n209), .C(n210), .D(n211), .Z(n207) );
  GTECH_OR_NOT U190 ( .A(n212), .B(n208), .Z(n211) );
  GTECH_XOR2 U191 ( .A(n213), .B(n152), .Z(n185) );
  GTECH_AND2 U192 ( .A(n214), .B(n215), .Z(n152) );
  GTECH_OR_NOT U193 ( .A(n216), .B(n217), .Z(n215) );
  GTECH_OAI21 U194 ( .A(n218), .B(n217), .C(n219), .Z(n214) );
  GTECH_OR_NOT U195 ( .A(n220), .B(I_a[7]), .Z(n213) );
  GTECH_NOT U196 ( .A(n161), .Z(n155) );
  GTECH_OAI2N2 U197 ( .A(n221), .B(n222), .C(n223), .D(n224), .Z(n161) );
  GTECH_OR_NOT U198 ( .A(n225), .B(n221), .Z(n224) );
  GTECH_XOR3 U199 ( .A(n221), .B(n225), .C(n226), .Z(N149) );
  GTECH_NOT U200 ( .A(n223), .Z(n226) );
  GTECH_XOR2 U201 ( .A(n227), .B(n188), .Z(n223) );
  GTECH_ADD_ABC U202 ( .A(n228), .B(n229), .C(n230), .COUT(n188) );
  GTECH_XOR3 U203 ( .A(n231), .B(n232), .C(n233), .Z(n229) );
  GTECH_OA21 U204 ( .A(n234), .B(n235), .C(n236), .Z(n228) );
  GTECH_XOR4 U205 ( .A(n193), .B(n205), .C(n203), .D(n191), .Z(n227) );
  GTECH_XOR3 U206 ( .A(n198), .B(n200), .C(n199), .Z(n191) );
  GTECH_OAI21 U207 ( .A(n237), .B(n238), .C(n239), .Z(n199) );
  GTECH_NOT U208 ( .A(n240), .Z(n200) );
  GTECH_OR_NOT U209 ( .A(n241), .B(I_b[7]), .Z(n240) );
  GTECH_NOT U210 ( .A(n196), .Z(n198) );
  GTECH_OR_NOT U211 ( .A(n202), .B(I_b[6]), .Z(n196) );
  GTECH_OR_NOT U212 ( .A(n179), .B(I_a[5]), .Z(n203) );
  GTECH_NOT U213 ( .A(I_b[4]), .Z(n179) );
  GTECH_OAI21 U214 ( .A(n233), .B(n242), .C(n243), .Z(n205) );
  GTECH_OAI21 U215 ( .A(n231), .B(n244), .C(n232), .Z(n243) );
  GTECH_NOT U216 ( .A(n242), .Z(n231) );
  GTECH_NOT U217 ( .A(n244), .Z(n233) );
  GTECH_NOT U218 ( .A(n245), .Z(n193) );
  GTECH_OR_NOT U219 ( .A(n178), .B(I_b[5]), .Z(n245) );
  GTECH_NOT U220 ( .A(n222), .Z(n225) );
  GTECH_XOR3 U221 ( .A(n212), .B(n208), .C(n210), .Z(n222) );
  GTECH_XOR3 U222 ( .A(n218), .B(n219), .C(n217), .Z(n210) );
  GTECH_OAI21 U223 ( .A(n246), .B(n247), .C(n248), .Z(n217) );
  GTECH_OAI21 U224 ( .A(n249), .B(n250), .C(n251), .Z(n248) );
  GTECH_NOT U225 ( .A(n250), .Z(n246) );
  GTECH_NOT U226 ( .A(n252), .Z(n219) );
  GTECH_OR_NOT U227 ( .A(n220), .B(I_a[6]), .Z(n252) );
  GTECH_NOT U228 ( .A(n216), .Z(n218) );
  GTECH_OR_NOT U229 ( .A(n253), .B(I_a[7]), .Z(n216) );
  GTECH_ADD_ABC U230 ( .A(n254), .B(n255), .C(n256), .COUT(n208) );
  GTECH_XOR2 U231 ( .A(n257), .B(n258), .Z(n255) );
  GTECH_AND2 U232 ( .A(I_a[7]), .B(I_b[1]), .Z(n258) );
  GTECH_NOT U233 ( .A(n209), .Z(n212) );
  GTECH_OR_NOT U234 ( .A(n257), .B(I_a[7]), .Z(n209) );
  GTECH_ADD_ABC U235 ( .A(n259), .B(n260), .C(n261), .COUT(n221) );
  GTECH_XOR3 U236 ( .A(n254), .B(n262), .C(n256), .Z(n260) );
  GTECH_NOT U237 ( .A(n263), .Z(n256) );
  GTECH_XOR2 U238 ( .A(n259), .B(n264), .Z(N148) );
  GTECH_XOR4 U239 ( .A(n262), .B(n263), .C(n261), .D(n254), .Z(n264) );
  GTECH_ADD_ABC U240 ( .A(n265), .B(n266), .C(n267), .COUT(n254) );
  GTECH_XOR3 U241 ( .A(n268), .B(n269), .C(n270), .Z(n266) );
  GTECH_XOR2 U242 ( .A(n271), .B(n272), .Z(n261) );
  GTECH_OA21 U243 ( .A(n234), .B(n235), .C(n236), .Z(n272) );
  GTECH_OAI21 U244 ( .A(n273), .B(n274), .C(n275), .Z(n236) );
  GTECH_NOT U245 ( .A(n234), .Z(n274) );
  GTECH_XOR4 U246 ( .A(n232), .B(n244), .C(n242), .D(n230), .Z(n271) );
  GTECH_XOR3 U247 ( .A(n276), .B(n277), .C(n239), .Z(n230) );
  GTECH_NAND3 U248 ( .A(I_b[6]), .B(I_a[1]), .C(n278), .Z(n239) );
  GTECH_NOT U249 ( .A(n238), .Z(n277) );
  GTECH_OR_NOT U250 ( .A(n279), .B(I_b[7]), .Z(n238) );
  GTECH_NOT U251 ( .A(n237), .Z(n276) );
  GTECH_OR_NOT U252 ( .A(n241), .B(I_b[6]), .Z(n237) );
  GTECH_OR_NOT U253 ( .A(n178), .B(I_b[4]), .Z(n242) );
  GTECH_OAI21 U254 ( .A(n280), .B(n281), .C(n282), .Z(n244) );
  GTECH_OAI21 U255 ( .A(n283), .B(n284), .C(n285), .Z(n282) );
  GTECH_NOT U256 ( .A(n284), .Z(n280) );
  GTECH_NOT U257 ( .A(n286), .Z(n232) );
  GTECH_OR_NOT U258 ( .A(n202), .B(I_b[5]), .Z(n286) );
  GTECH_XOR3 U259 ( .A(n249), .B(n251), .C(n250), .Z(n263) );
  GTECH_OAI21 U260 ( .A(n287), .B(n288), .C(n289), .Z(n250) );
  GTECH_OAI21 U261 ( .A(n290), .B(n291), .C(n292), .Z(n289) );
  GTECH_NOT U262 ( .A(n291), .Z(n287) );
  GTECH_NOT U263 ( .A(n293), .Z(n251) );
  GTECH_OR_NOT U264 ( .A(n220), .B(I_a[5]), .Z(n293) );
  GTECH_NOT U265 ( .A(I_b[3]), .Z(n220) );
  GTECH_NOT U266 ( .A(n247), .Z(n249) );
  GTECH_OR_NOT U267 ( .A(n253), .B(I_a[6]), .Z(n247) );
  GTECH_XOR2 U268 ( .A(n294), .B(n257), .Z(n262) );
  GTECH_OA21 U269 ( .A(n270), .B(n295), .C(n296), .Z(n257) );
  GTECH_OAI21 U270 ( .A(n268), .B(n297), .C(n269), .Z(n296) );
  GTECH_NOT U271 ( .A(n297), .Z(n270) );
  GTECH_AND2 U272 ( .A(I_b[1]), .B(I_a[7]), .Z(n294) );
  GTECH_ADD_ABC U273 ( .A(n298), .B(n299), .C(n300), .COUT(n259) );
  GTECH_NOT U274 ( .A(n301), .Z(n300) );
  GTECH_XOR3 U275 ( .A(n265), .B(n302), .C(n267), .Z(n299) );
  GTECH_NOT U276 ( .A(n303), .Z(n267) );
  GTECH_NOT U277 ( .A(n304), .Z(n302) );
  GTECH_XOR2 U278 ( .A(n305), .B(n298), .Z(N147) );
  GTECH_ADD_ABC U279 ( .A(n306), .B(n307), .C(n308), .COUT(n298) );
  GTECH_XOR3 U280 ( .A(n309), .B(n310), .C(n311), .Z(n307) );
  GTECH_OA21 U281 ( .A(n312), .B(n313), .C(n314), .Z(n306) );
  GTECH_XOR4 U282 ( .A(n303), .B(n265), .C(n304), .D(n301), .Z(n305) );
  GTECH_XOR3 U283 ( .A(n275), .B(n235), .C(n234), .Z(n301) );
  GTECH_XOR2 U284 ( .A(n315), .B(n278), .Z(n234) );
  GTECH_NOT U285 ( .A(n316), .Z(n278) );
  GTECH_OR_NOT U286 ( .A(n317), .B(I_b[7]), .Z(n316) );
  GTECH_OR_NOT U287 ( .A(n279), .B(I_b[6]), .Z(n315) );
  GTECH_NOT U288 ( .A(n273), .Z(n235) );
  GTECH_XOR3 U289 ( .A(n283), .B(n285), .C(n284), .Z(n273) );
  GTECH_OAI21 U290 ( .A(n318), .B(n319), .C(n320), .Z(n284) );
  GTECH_NOT U291 ( .A(n321), .Z(n285) );
  GTECH_OR_NOT U292 ( .A(n241), .B(I_b[5]), .Z(n321) );
  GTECH_NOT U293 ( .A(n281), .Z(n283) );
  GTECH_OR_NOT U294 ( .A(n202), .B(I_b[4]), .Z(n281) );
  GTECH_NOT U295 ( .A(n322), .Z(n275) );
  GTECH_NAND3 U296 ( .A(I_a[0]), .B(n323), .C(I_b[6]), .Z(n322) );
  GTECH_NOT U297 ( .A(n324), .Z(n323) );
  GTECH_XOR3 U298 ( .A(n268), .B(n269), .C(n297), .Z(n304) );
  GTECH_OAI21 U299 ( .A(n325), .B(n326), .C(n327), .Z(n297) );
  GTECH_OAI21 U300 ( .A(n328), .B(n329), .C(n330), .Z(n327) );
  GTECH_NOT U301 ( .A(n331), .Z(n269) );
  GTECH_OR_NOT U302 ( .A(n332), .B(I_a[6]), .Z(n331) );
  GTECH_NOT U303 ( .A(n295), .Z(n268) );
  GTECH_OR_NOT U304 ( .A(n333), .B(I_a[7]), .Z(n295) );
  GTECH_ADD_ABC U305 ( .A(n309), .B(n334), .C(n311), .COUT(n265) );
  GTECH_NOT U306 ( .A(n335), .Z(n311) );
  GTECH_XOR3 U307 ( .A(n328), .B(n330), .C(n325), .Z(n334) );
  GTECH_NOT U308 ( .A(n329), .Z(n325) );
  GTECH_XOR3 U309 ( .A(n290), .B(n292), .C(n291), .Z(n303) );
  GTECH_OAI21 U310 ( .A(n336), .B(n337), .C(n338), .Z(n291) );
  GTECH_OAI21 U311 ( .A(n339), .B(n340), .C(n341), .Z(n338) );
  GTECH_NOT U312 ( .A(n340), .Z(n336) );
  GTECH_NOT U313 ( .A(n342), .Z(n292) );
  GTECH_OR_NOT U314 ( .A(n178), .B(I_b[3]), .Z(n342) );
  GTECH_NOT U315 ( .A(n288), .Z(n290) );
  GTECH_OR_NOT U316 ( .A(n253), .B(I_a[5]), .Z(n288) );
  GTECH_NOT U317 ( .A(I_b[2]), .Z(n253) );
  GTECH_XOR2 U318 ( .A(n343), .B(n344), .Z(N146) );
  GTECH_XOR4 U319 ( .A(n310), .B(n335), .C(n308), .D(n309), .Z(n344) );
  GTECH_ADD_ABC U320 ( .A(n345), .B(n346), .C(n347), .COUT(n309) );
  GTECH_NOT U321 ( .A(n348), .Z(n347) );
  GTECH_XOR3 U322 ( .A(n349), .B(n350), .C(n351), .Z(n346) );
  GTECH_XOR2 U323 ( .A(n324), .B(n352), .Z(n308) );
  GTECH_AND2 U324 ( .A(I_b[6]), .B(I_a[0]), .Z(n352) );
  GTECH_XOR3 U325 ( .A(n353), .B(n354), .C(n320), .Z(n324) );
  GTECH_NAND3 U326 ( .A(I_b[4]), .B(I_a[1]), .C(n355), .Z(n320) );
  GTECH_NOT U327 ( .A(n319), .Z(n354) );
  GTECH_OR_NOT U328 ( .A(n279), .B(I_b[5]), .Z(n319) );
  GTECH_NOT U329 ( .A(n318), .Z(n353) );
  GTECH_OR_NOT U330 ( .A(n241), .B(I_b[4]), .Z(n318) );
  GTECH_XOR3 U331 ( .A(n339), .B(n341), .C(n340), .Z(n335) );
  GTECH_OAI21 U332 ( .A(n356), .B(n357), .C(n358), .Z(n340) );
  GTECH_OAI21 U333 ( .A(n359), .B(n360), .C(n361), .Z(n358) );
  GTECH_NOT U334 ( .A(n360), .Z(n356) );
  GTECH_NOT U335 ( .A(n362), .Z(n341) );
  GTECH_OR_NOT U336 ( .A(n202), .B(I_b[3]), .Z(n362) );
  GTECH_NOT U337 ( .A(n337), .Z(n339) );
  GTECH_OR_NOT U338 ( .A(n178), .B(I_b[2]), .Z(n337) );
  GTECH_NOT U339 ( .A(I_a[4]), .Z(n178) );
  GTECH_NOT U340 ( .A(n363), .Z(n310) );
  GTECH_XOR3 U341 ( .A(n328), .B(n330), .C(n329), .Z(n363) );
  GTECH_OAI21 U342 ( .A(n351), .B(n364), .C(n365), .Z(n329) );
  GTECH_OAI21 U343 ( .A(n349), .B(n366), .C(n350), .Z(n365) );
  GTECH_NOT U344 ( .A(n364), .Z(n349) );
  GTECH_NOT U345 ( .A(n366), .Z(n351) );
  GTECH_NOT U346 ( .A(n367), .Z(n330) );
  GTECH_OR_NOT U347 ( .A(n332), .B(I_a[5]), .Z(n367) );
  GTECH_NOT U348 ( .A(n326), .Z(n328) );
  GTECH_OR_NOT U349 ( .A(n333), .B(I_a[6]), .Z(n326) );
  GTECH_OA21 U350 ( .A(n312), .B(n313), .C(n314), .Z(n343) );
  GTECH_OAI21 U351 ( .A(n368), .B(n369), .C(n370), .Z(n314) );
  GTECH_NOT U352 ( .A(n312), .Z(n369) );
  GTECH_XOR3 U353 ( .A(n370), .B(n313), .C(n312), .Z(N145) );
  GTECH_XOR2 U354 ( .A(n371), .B(n355), .Z(n312) );
  GTECH_NOT U355 ( .A(n372), .Z(n355) );
  GTECH_OR_NOT U356 ( .A(n317), .B(I_b[5]), .Z(n372) );
  GTECH_OR_NOT U357 ( .A(n279), .B(I_b[4]), .Z(n371) );
  GTECH_NOT U358 ( .A(n368), .Z(n313) );
  GTECH_XOR2 U359 ( .A(n373), .B(n345), .Z(n368) );
  GTECH_ADD_ABC U360 ( .A(n374), .B(n375), .C(n376), .COUT(n345) );
  GTECH_XOR3 U361 ( .A(n377), .B(n378), .C(n379), .Z(n375) );
  GTECH_OA21 U362 ( .A(n380), .B(n381), .C(n382), .Z(n374) );
  GTECH_XOR4 U363 ( .A(n350), .B(n366), .C(n364), .D(n348), .Z(n373) );
  GTECH_XOR3 U364 ( .A(n359), .B(n361), .C(n360), .Z(n348) );
  GTECH_OAI21 U365 ( .A(n383), .B(n384), .C(n385), .Z(n360) );
  GTECH_NOT U366 ( .A(n386), .Z(n361) );
  GTECH_OR_NOT U367 ( .A(n241), .B(I_b[3]), .Z(n386) );
  GTECH_NOT U368 ( .A(n357), .Z(n359) );
  GTECH_OR_NOT U369 ( .A(n202), .B(I_b[2]), .Z(n357) );
  GTECH_OR_NOT U370 ( .A(n333), .B(I_a[5]), .Z(n364) );
  GTECH_OAI21 U371 ( .A(n379), .B(n387), .C(n388), .Z(n366) );
  GTECH_OAI21 U372 ( .A(n377), .B(n389), .C(n378), .Z(n388) );
  GTECH_NOT U373 ( .A(n389), .Z(n379) );
  GTECH_NOT U374 ( .A(n390), .Z(n350) );
  GTECH_OR_NOT U375 ( .A(n332), .B(I_a[4]), .Z(n390) );
  GTECH_NOT U376 ( .A(n391), .Z(n370) );
  GTECH_NAND3 U377 ( .A(I_a[0]), .B(n392), .C(I_b[4]), .Z(n391) );
  GTECH_XOR2 U378 ( .A(n393), .B(n392), .Z(N144) );
  GTECH_XOR2 U379 ( .A(n394), .B(n395), .Z(n392) );
  GTECH_XOR4 U380 ( .A(n378), .B(n389), .C(n376), .D(n377), .Z(n395) );
  GTECH_NOT U381 ( .A(n387), .Z(n377) );
  GTECH_OR_NOT U382 ( .A(n333), .B(I_a[4]), .Z(n387) );
  GTECH_NOT U383 ( .A(I_b[0]), .Z(n333) );
  GTECH_XOR3 U384 ( .A(n396), .B(n397), .C(n385), .Z(n376) );
  GTECH_NAND3 U385 ( .A(I_b[2]), .B(I_a[1]), .C(n398), .Z(n385) );
  GTECH_NOT U386 ( .A(n384), .Z(n397) );
  GTECH_OR_NOT U387 ( .A(n279), .B(I_b[3]), .Z(n384) );
  GTECH_NOT U388 ( .A(n383), .Z(n396) );
  GTECH_OR_NOT U389 ( .A(n241), .B(I_b[2]), .Z(n383) );
  GTECH_OAI21 U390 ( .A(n399), .B(n400), .C(n401), .Z(n389) );
  GTECH_OAI21 U391 ( .A(n402), .B(n403), .C(n404), .Z(n401) );
  GTECH_NOT U392 ( .A(n403), .Z(n399) );
  GTECH_NOT U393 ( .A(n405), .Z(n378) );
  GTECH_OR_NOT U394 ( .A(n332), .B(I_a[3]), .Z(n405) );
  GTECH_OA21 U395 ( .A(n380), .B(n381), .C(n382), .Z(n394) );
  GTECH_OAI21 U396 ( .A(n406), .B(n407), .C(n408), .Z(n382) );
  GTECH_NOT U397 ( .A(n380), .Z(n407) );
  GTECH_AND2 U398 ( .A(I_b[4]), .B(I_a[0]), .Z(n393) );
  GTECH_XOR3 U399 ( .A(n408), .B(n381), .C(n380), .Z(N143) );
  GTECH_XOR2 U400 ( .A(n409), .B(n398), .Z(n380) );
  GTECH_NOT U401 ( .A(n410), .Z(n398) );
  GTECH_OR_NOT U402 ( .A(n317), .B(I_b[3]), .Z(n410) );
  GTECH_NOT U403 ( .A(I_a[0]), .Z(n317) );
  GTECH_OR_NOT U404 ( .A(n279), .B(I_b[2]), .Z(n409) );
  GTECH_NOT U405 ( .A(I_a[1]), .Z(n279) );
  GTECH_NOT U406 ( .A(n406), .Z(n381) );
  GTECH_XOR3 U407 ( .A(n402), .B(n404), .C(n403), .Z(n406) );
  GTECH_OAI21 U408 ( .A(n411), .B(n412), .C(n413), .Z(n403) );
  GTECH_NOT U409 ( .A(n414), .Z(n404) );
  GTECH_OR_NOT U410 ( .A(n241), .B(I_b[1]), .Z(n414) );
  GTECH_NOT U411 ( .A(n400), .Z(n402) );
  GTECH_OR_NOT U412 ( .A(n202), .B(I_b[0]), .Z(n400) );
  GTECH_NOT U413 ( .A(I_a[3]), .Z(n202) );
  GTECH_NOT U414 ( .A(n415), .Z(n408) );
  GTECH_NAND3 U415 ( .A(I_a[0]), .B(n416), .C(I_b[2]), .Z(n415) );
  GTECH_XOR2 U416 ( .A(n417), .B(n416), .Z(N142) );
  GTECH_NOT U417 ( .A(n418), .Z(n416) );
  GTECH_XOR3 U418 ( .A(n419), .B(n420), .C(n413), .Z(n418) );
  GTECH_NAND3 U419 ( .A(n421), .B(I_b[0]), .C(I_a[1]), .Z(n413) );
  GTECH_NOT U420 ( .A(n411), .Z(n420) );
  GTECH_OR_NOT U421 ( .A(n332), .B(I_a[1]), .Z(n411) );
  GTECH_NOT U422 ( .A(n412), .Z(n419) );
  GTECH_OR_NOT U423 ( .A(n241), .B(I_b[0]), .Z(n412) );
  GTECH_NOT U424 ( .A(I_a[2]), .Z(n241) );
  GTECH_AND2 U425 ( .A(I_b[2]), .B(I_a[0]), .Z(n417) );
  GTECH_XOR2 U426 ( .A(n421), .B(n422), .Z(N141) );
  GTECH_AND2 U427 ( .A(I_a[1]), .B(I_b[0]), .Z(n422) );
  GTECH_NOT U428 ( .A(n423), .Z(n421) );
  GTECH_OR_NOT U429 ( .A(n332), .B(I_a[0]), .Z(n423) );
  GTECH_NOT U430 ( .A(I_b[1]), .Z(n332) );
  GTECH_AND2 U431 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

