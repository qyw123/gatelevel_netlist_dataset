
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NAND2 U83 ( .A(n93), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI21 U86 ( .A(n98), .B(n99), .C(n100), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_NAND2 U88 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U89 ( .A(n104), .Z(n84) );
  GTECH_NAND2 U90 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_XOR2 U91 ( .A(n106), .B(n105), .Z(N153) );
  GTECH_NOT U92 ( .A(n107), .Z(n105) );
  GTECH_XNOR3 U93 ( .A(n108), .B(n93), .C(n109), .Z(n107) );
  GTECH_NOT U94 ( .A(n95), .Z(n109) );
  GTECH_XNOR3 U95 ( .A(n101), .B(n103), .C(n98), .Z(n95) );
  GTECH_NOT U96 ( .A(n102), .Z(n98) );
  GTECH_OAI21 U97 ( .A(n110), .B(n111), .C(n112), .Z(n102) );
  GTECH_OAI21 U98 ( .A(n113), .B(n114), .C(n115), .Z(n112) );
  GTECH_NOT U99 ( .A(n116), .Z(n103) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n116) );
  GTECH_NOT U101 ( .A(n99), .Z(n101) );
  GTECH_NAND2 U102 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U103 ( .A(n117), .B(n118), .C(n119), .COUT(n93) );
  GTECH_NOT U104 ( .A(n120), .Z(n119) );
  GTECH_XOR2 U105 ( .A(n121), .B(n122), .Z(n118) );
  GTECH_AND2 U106 ( .A(I_a[7]), .B(I_b[5]), .Z(n122) );
  GTECH_NOT U107 ( .A(n94), .Z(n108) );
  GTECH_NAND2 U108 ( .A(I_a[7]), .B(n123), .Z(n94) );
  GTECH_NOT U109 ( .A(n124), .Z(n106) );
  GTECH_NAND2 U110 ( .A(n125), .B(n126), .Z(n124) );
  GTECH_NOT U111 ( .A(n127), .Z(n126) );
  GTECH_XOR2 U112 ( .A(n127), .B(n128), .Z(N152) );
  GTECH_NOT U113 ( .A(n125), .Z(n128) );
  GTECH_XOR4 U114 ( .A(n129), .B(n121), .C(n120), .D(n117), .Z(n125) );
  GTECH_ADD_ABC U115 ( .A(n130), .B(n131), .C(n132), .COUT(n117) );
  GTECH_XNOR3 U116 ( .A(n133), .B(n134), .C(n135), .Z(n131) );
  GTECH_XNOR3 U117 ( .A(n113), .B(n115), .C(n110), .Z(n120) );
  GTECH_NOT U118 ( .A(n114), .Z(n110) );
  GTECH_OAI21 U119 ( .A(n136), .B(n137), .C(n138), .Z(n114) );
  GTECH_OAI21 U120 ( .A(n139), .B(n140), .C(n141), .Z(n138) );
  GTECH_NOT U121 ( .A(n142), .Z(n115) );
  GTECH_NAND2 U122 ( .A(I_b[7]), .B(I_a[5]), .Z(n142) );
  GTECH_NOT U123 ( .A(n111), .Z(n113) );
  GTECH_NAND2 U124 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_NOT U125 ( .A(n123), .Z(n121) );
  GTECH_OAI21 U126 ( .A(n143), .B(n144), .C(n145), .Z(n123) );
  GTECH_OAI21 U127 ( .A(n133), .B(n135), .C(n134), .Z(n145) );
  GTECH_AND2 U128 ( .A(I_a[7]), .B(I_b[5]), .Z(n129) );
  GTECH_ADD_ABC U129 ( .A(n146), .B(n147), .C(n148), .COUT(n127) );
  GTECH_AOI2N2 U130 ( .A(n149), .B(n150), .C(n151), .D(n152), .Z(n148) );
  GTECH_NAND2 U131 ( .A(n152), .B(n151), .Z(n149) );
  GTECH_OA22 U132 ( .A(n153), .B(n154), .C(n155), .D(n156), .Z(n147) );
  GTECH_XNOR3 U133 ( .A(n157), .B(n146), .C(n158), .Z(N151) );
  GTECH_AOI2N2 U134 ( .A(n150), .B(n159), .C(n152), .D(n151), .Z(n158) );
  GTECH_OR_NOT U135 ( .A(n160), .B(n151), .Z(n159) );
  GTECH_XOR2 U136 ( .A(n130), .B(n161), .Z(n146) );
  GTECH_XOR4 U137 ( .A(n134), .B(n143), .C(n132), .D(n133), .Z(n161) );
  GTECH_NOT U138 ( .A(n144), .Z(n133) );
  GTECH_NAND2 U139 ( .A(I_a[7]), .B(I_b[4]), .Z(n144) );
  GTECH_NOT U140 ( .A(n162), .Z(n132) );
  GTECH_XNOR3 U141 ( .A(n139), .B(n141), .C(n136), .Z(n162) );
  GTECH_NOT U142 ( .A(n140), .Z(n136) );
  GTECH_OAI21 U143 ( .A(n163), .B(n164), .C(n165), .Z(n140) );
  GTECH_OAI21 U144 ( .A(n166), .B(n167), .C(n168), .Z(n165) );
  GTECH_NOT U145 ( .A(n169), .Z(n141) );
  GTECH_NAND2 U146 ( .A(I_b[7]), .B(I_a[4]), .Z(n169) );
  GTECH_NOT U147 ( .A(n137), .Z(n139) );
  GTECH_NAND2 U148 ( .A(I_b[6]), .B(I_a[5]), .Z(n137) );
  GTECH_NOT U149 ( .A(n135), .Z(n143) );
  GTECH_OAI21 U150 ( .A(n170), .B(n171), .C(n172), .Z(n135) );
  GTECH_OAI21 U151 ( .A(n173), .B(n174), .C(n175), .Z(n172) );
  GTECH_NOT U152 ( .A(n176), .Z(n134) );
  GTECH_NAND2 U153 ( .A(I_a[6]), .B(I_b[5]), .Z(n176) );
  GTECH_ADD_ABC U154 ( .A(n177), .B(n178), .C(n179), .COUT(n130) );
  GTECH_NOT U155 ( .A(n180), .Z(n179) );
  GTECH_XNOR3 U156 ( .A(n173), .B(n175), .C(n174), .Z(n178) );
  GTECH_OA22 U157 ( .A(n156), .B(n155), .C(n154), .D(n153), .Z(n157) );
  GTECH_NOT U158 ( .A(n181), .Z(n153) );
  GTECH_NOT U159 ( .A(I_a[7]), .Z(n155) );
  GTECH_XNOR3 U160 ( .A(n152), .B(n182), .C(n150), .Z(N150) );
  GTECH_XOR2 U161 ( .A(n183), .B(n177), .Z(n150) );
  GTECH_ADD_ABC U162 ( .A(n184), .B(n185), .C(n186), .COUT(n177) );
  GTECH_NOT U163 ( .A(n187), .Z(n186) );
  GTECH_XNOR3 U164 ( .A(n188), .B(n189), .C(n190), .Z(n185) );
  GTECH_XOR4 U165 ( .A(n175), .B(n170), .C(n180), .D(n173), .Z(n183) );
  GTECH_NOT U166 ( .A(n171), .Z(n173) );
  GTECH_NAND2 U167 ( .A(I_a[6]), .B(I_b[4]), .Z(n171) );
  GTECH_XNOR3 U168 ( .A(n166), .B(n168), .C(n163), .Z(n180) );
  GTECH_NOT U169 ( .A(n167), .Z(n163) );
  GTECH_OAI21 U170 ( .A(n191), .B(n192), .C(n193), .Z(n167) );
  GTECH_OAI21 U171 ( .A(n194), .B(n195), .C(n196), .Z(n193) );
  GTECH_NOT U172 ( .A(n197), .Z(n168) );
  GTECH_NAND2 U173 ( .A(I_b[7]), .B(I_a[3]), .Z(n197) );
  GTECH_NOT U174 ( .A(n164), .Z(n166) );
  GTECH_NAND2 U175 ( .A(I_b[6]), .B(I_a[4]), .Z(n164) );
  GTECH_NOT U176 ( .A(n174), .Z(n170) );
  GTECH_OAI21 U177 ( .A(n198), .B(n199), .C(n200), .Z(n174) );
  GTECH_OAI21 U178 ( .A(n188), .B(n190), .C(n189), .Z(n200) );
  GTECH_NOT U179 ( .A(n201), .Z(n175) );
  GTECH_NAND2 U180 ( .A(I_a[5]), .B(I_b[5]), .Z(n201) );
  GTECH_NOT U181 ( .A(n151), .Z(n182) );
  GTECH_XOR2 U182 ( .A(n181), .B(n154), .Z(n151) );
  GTECH_AOI2N2 U183 ( .A(n202), .B(n203), .C(n204), .D(n205), .Z(n154) );
  GTECH_NAND2 U184 ( .A(n204), .B(n205), .Z(n203) );
  GTECH_XOR2 U185 ( .A(n206), .B(n156), .Z(n181) );
  GTECH_OA22 U186 ( .A(n207), .B(n208), .C(n209), .D(n210), .Z(n156) );
  GTECH_AND_NOT U187 ( .A(n208), .B(n211), .Z(n209) );
  GTECH_NAND2 U188 ( .A(I_a[7]), .B(I_b[3]), .Z(n206) );
  GTECH_NOT U189 ( .A(n160), .Z(n152) );
  GTECH_OAI2N2 U190 ( .A(n212), .B(n213), .C(n214), .D(n215), .Z(n160) );
  GTECH_NAND2 U191 ( .A(n212), .B(n213), .Z(n215) );
  GTECH_XNOR3 U192 ( .A(n212), .B(n216), .C(n214), .Z(N149) );
  GTECH_XOR2 U193 ( .A(n217), .B(n184), .Z(n214) );
  GTECH_ADD_ABC U194 ( .A(n218), .B(n219), .C(n220), .COUT(n184) );
  GTECH_XNOR3 U195 ( .A(n221), .B(n222), .C(n223), .Z(n219) );
  GTECH_OA22 U196 ( .A(n224), .B(n225), .C(n226), .D(n227), .Z(n218) );
  GTECH_AND2 U197 ( .A(n226), .B(n227), .Z(n224) );
  GTECH_XOR4 U198 ( .A(n189), .B(n198), .C(n187), .D(n188), .Z(n217) );
  GTECH_NOT U199 ( .A(n199), .Z(n188) );
  GTECH_NAND2 U200 ( .A(I_a[5]), .B(I_b[4]), .Z(n199) );
  GTECH_XNOR3 U201 ( .A(n194), .B(n196), .C(n191), .Z(n187) );
  GTECH_NOT U202 ( .A(n195), .Z(n191) );
  GTECH_OAI21 U203 ( .A(n228), .B(n229), .C(n230), .Z(n195) );
  GTECH_NOT U204 ( .A(n231), .Z(n196) );
  GTECH_NAND2 U205 ( .A(I_b[7]), .B(I_a[2]), .Z(n231) );
  GTECH_NOT U206 ( .A(n192), .Z(n194) );
  GTECH_NAND2 U207 ( .A(I_b[6]), .B(I_a[3]), .Z(n192) );
  GTECH_NOT U208 ( .A(n190), .Z(n198) );
  GTECH_OAI21 U209 ( .A(n232), .B(n233), .C(n234), .Z(n190) );
  GTECH_OAI21 U210 ( .A(n221), .B(n223), .C(n222), .Z(n234) );
  GTECH_NOT U211 ( .A(n235), .Z(n189) );
  GTECH_NAND2 U212 ( .A(I_b[5]), .B(I_a[4]), .Z(n235) );
  GTECH_NOT U213 ( .A(n213), .Z(n216) );
  GTECH_XNOR3 U214 ( .A(n236), .B(n204), .C(n237), .Z(n213) );
  GTECH_NOT U215 ( .A(n202), .Z(n237) );
  GTECH_XNOR3 U216 ( .A(n238), .B(n239), .C(n207), .Z(n202) );
  GTECH_NOT U217 ( .A(n211), .Z(n207) );
  GTECH_OAI21 U218 ( .A(n240), .B(n241), .C(n242), .Z(n211) );
  GTECH_OAI21 U219 ( .A(n243), .B(n244), .C(n245), .Z(n242) );
  GTECH_NOT U220 ( .A(n210), .Z(n239) );
  GTECH_NAND2 U221 ( .A(I_a[6]), .B(I_b[3]), .Z(n210) );
  GTECH_NOT U222 ( .A(n208), .Z(n238) );
  GTECH_NAND2 U223 ( .A(I_a[7]), .B(I_b[2]), .Z(n208) );
  GTECH_ADD_ABC U224 ( .A(n246), .B(n247), .C(n248), .COUT(n204) );
  GTECH_NOT U225 ( .A(n249), .Z(n248) );
  GTECH_XOR2 U226 ( .A(n250), .B(n251), .Z(n247) );
  GTECH_AND2 U227 ( .A(I_a[7]), .B(I_b[1]), .Z(n251) );
  GTECH_NOT U228 ( .A(n205), .Z(n236) );
  GTECH_NAND2 U229 ( .A(I_a[7]), .B(n252), .Z(n205) );
  GTECH_ADD_ABC U230 ( .A(n253), .B(n254), .C(n255), .COUT(n212) );
  GTECH_XNOR3 U231 ( .A(n246), .B(n256), .C(n249), .Z(n254) );
  GTECH_XOR2 U232 ( .A(n257), .B(n253), .Z(N148) );
  GTECH_ADD_ABC U233 ( .A(n258), .B(n259), .C(n260), .COUT(n253) );
  GTECH_NOT U234 ( .A(n261), .Z(n260) );
  GTECH_XNOR3 U235 ( .A(n262), .B(n263), .C(n264), .Z(n259) );
  GTECH_XOR4 U236 ( .A(n256), .B(n246), .C(n249), .D(n255), .Z(n257) );
  GTECH_XOR2 U237 ( .A(n265), .B(n266), .Z(n255) );
  GTECH_XOR4 U238 ( .A(n222), .B(n232), .C(n220), .D(n221), .Z(n266) );
  GTECH_NOT U239 ( .A(n233), .Z(n221) );
  GTECH_NAND2 U240 ( .A(I_b[4]), .B(I_a[4]), .Z(n233) );
  GTECH_XNOR3 U241 ( .A(n267), .B(n268), .C(n269), .Z(n220) );
  GTECH_NOT U242 ( .A(n230), .Z(n269) );
  GTECH_NAND3 U243 ( .A(I_b[6]), .B(I_a[1]), .C(n270), .Z(n230) );
  GTECH_NOT U244 ( .A(n229), .Z(n268) );
  GTECH_NAND2 U245 ( .A(I_b[7]), .B(I_a[1]), .Z(n229) );
  GTECH_NOT U246 ( .A(n228), .Z(n267) );
  GTECH_NAND2 U247 ( .A(I_b[6]), .B(I_a[2]), .Z(n228) );
  GTECH_NOT U248 ( .A(n223), .Z(n232) );
  GTECH_OAI21 U249 ( .A(n271), .B(n272), .C(n273), .Z(n223) );
  GTECH_OAI21 U250 ( .A(n274), .B(n275), .C(n276), .Z(n273) );
  GTECH_NOT U251 ( .A(n277), .Z(n222) );
  GTECH_NAND2 U252 ( .A(I_b[5]), .B(I_a[3]), .Z(n277) );
  GTECH_OA22 U253 ( .A(n226), .B(n227), .C(n278), .D(n225), .Z(n265) );
  GTECH_AND_NOT U254 ( .A(n226), .B(n279), .Z(n278) );
  GTECH_XNOR3 U255 ( .A(n243), .B(n245), .C(n240), .Z(n249) );
  GTECH_NOT U256 ( .A(n244), .Z(n240) );
  GTECH_OAI21 U257 ( .A(n280), .B(n281), .C(n282), .Z(n244) );
  GTECH_OAI21 U258 ( .A(n283), .B(n284), .C(n285), .Z(n282) );
  GTECH_NOT U259 ( .A(n286), .Z(n245) );
  GTECH_NAND2 U260 ( .A(I_a[5]), .B(I_b[3]), .Z(n286) );
  GTECH_NOT U261 ( .A(n241), .Z(n243) );
  GTECH_NAND2 U262 ( .A(I_a[6]), .B(I_b[2]), .Z(n241) );
  GTECH_ADD_ABC U263 ( .A(n262), .B(n287), .C(n288), .COUT(n246) );
  GTECH_XNOR3 U264 ( .A(n289), .B(n290), .C(n291), .Z(n287) );
  GTECH_XOR2 U265 ( .A(n292), .B(n250), .Z(n256) );
  GTECH_NOT U266 ( .A(n252), .Z(n250) );
  GTECH_OAI21 U267 ( .A(n293), .B(n294), .C(n295), .Z(n252) );
  GTECH_OAI21 U268 ( .A(n289), .B(n291), .C(n290), .Z(n295) );
  GTECH_AND2 U269 ( .A(I_a[7]), .B(I_b[1]), .Z(n292) );
  GTECH_XOR2 U270 ( .A(n296), .B(n258), .Z(N147) );
  GTECH_ADD_ABC U271 ( .A(n297), .B(n298), .C(n299), .COUT(n258) );
  GTECH_XNOR3 U272 ( .A(n300), .B(n301), .C(n302), .Z(n298) );
  GTECH_OA22 U273 ( .A(n303), .B(n304), .C(n305), .D(n306), .Z(n297) );
  GTECH_AND2 U274 ( .A(n305), .B(n306), .Z(n303) );
  GTECH_XOR4 U275 ( .A(n263), .B(n288), .C(n261), .D(n262), .Z(n296) );
  GTECH_ADD_ABC U276 ( .A(n300), .B(n307), .C(n308), .COUT(n262) );
  GTECH_NOT U277 ( .A(n302), .Z(n308) );
  GTECH_XNOR3 U278 ( .A(n309), .B(n310), .C(n311), .Z(n307) );
  GTECH_XNOR3 U279 ( .A(n312), .B(n227), .C(n313), .Z(n261) );
  GTECH_NOT U280 ( .A(n226), .Z(n313) );
  GTECH_XOR2 U281 ( .A(n314), .B(n270), .Z(n226) );
  GTECH_NOT U282 ( .A(n315), .Z(n270) );
  GTECH_NAND2 U283 ( .A(I_b[7]), .B(I_a[0]), .Z(n315) );
  GTECH_NAND2 U284 ( .A(I_b[6]), .B(I_a[1]), .Z(n314) );
  GTECH_NOT U285 ( .A(n279), .Z(n227) );
  GTECH_XNOR3 U286 ( .A(n274), .B(n276), .C(n271), .Z(n279) );
  GTECH_NOT U287 ( .A(n275), .Z(n271) );
  GTECH_OAI21 U288 ( .A(n316), .B(n317), .C(n318), .Z(n275) );
  GTECH_NOT U289 ( .A(n319), .Z(n276) );
  GTECH_NAND2 U290 ( .A(I_b[5]), .B(I_a[2]), .Z(n319) );
  GTECH_NOT U291 ( .A(n272), .Z(n274) );
  GTECH_NAND2 U292 ( .A(I_b[4]), .B(I_a[3]), .Z(n272) );
  GTECH_NOT U293 ( .A(n225), .Z(n312) );
  GTECH_NAND3 U294 ( .A(I_a[0]), .B(n320), .C(I_b[6]), .Z(n225) );
  GTECH_NOT U295 ( .A(n321), .Z(n320) );
  GTECH_NOT U296 ( .A(n264), .Z(n288) );
  GTECH_XNOR3 U297 ( .A(n283), .B(n285), .C(n280), .Z(n264) );
  GTECH_NOT U298 ( .A(n284), .Z(n280) );
  GTECH_OAI21 U299 ( .A(n322), .B(n323), .C(n324), .Z(n284) );
  GTECH_OAI21 U300 ( .A(n325), .B(n326), .C(n327), .Z(n324) );
  GTECH_NOT U301 ( .A(n328), .Z(n285) );
  GTECH_NAND2 U302 ( .A(I_b[3]), .B(I_a[4]), .Z(n328) );
  GTECH_NOT U303 ( .A(n281), .Z(n283) );
  GTECH_NAND2 U304 ( .A(I_a[5]), .B(I_b[2]), .Z(n281) );
  GTECH_NOT U305 ( .A(n329), .Z(n263) );
  GTECH_XNOR3 U306 ( .A(n289), .B(n290), .C(n293), .Z(n329) );
  GTECH_NOT U307 ( .A(n291), .Z(n293) );
  GTECH_OAI21 U308 ( .A(n330), .B(n331), .C(n332), .Z(n291) );
  GTECH_OAI21 U309 ( .A(n309), .B(n311), .C(n310), .Z(n332) );
  GTECH_NOT U310 ( .A(n333), .Z(n290) );
  GTECH_NAND2 U311 ( .A(I_a[6]), .B(I_b[1]), .Z(n333) );
  GTECH_NOT U312 ( .A(n294), .Z(n289) );
  GTECH_NAND2 U313 ( .A(I_a[7]), .B(I_b[0]), .Z(n294) );
  GTECH_XOR2 U314 ( .A(n334), .B(n335), .Z(N146) );
  GTECH_OA22 U315 ( .A(n305), .B(n306), .C(n336), .D(n304), .Z(n335) );
  GTECH_AND_NOT U316 ( .A(n305), .B(n337), .Z(n336) );
  GTECH_XOR4 U317 ( .A(n301), .B(n300), .C(n302), .D(n299), .Z(n334) );
  GTECH_XOR2 U318 ( .A(n321), .B(n338), .Z(n299) );
  GTECH_AND2 U319 ( .A(I_b[6]), .B(I_a[0]), .Z(n338) );
  GTECH_XNOR3 U320 ( .A(n339), .B(n340), .C(n341), .Z(n321) );
  GTECH_NOT U321 ( .A(n318), .Z(n341) );
  GTECH_NAND3 U322 ( .A(I_b[4]), .B(I_a[1]), .C(n342), .Z(n318) );
  GTECH_NOT U323 ( .A(n317), .Z(n340) );
  GTECH_NAND2 U324 ( .A(I_b[5]), .B(I_a[1]), .Z(n317) );
  GTECH_NOT U325 ( .A(n316), .Z(n339) );
  GTECH_NAND2 U326 ( .A(I_b[4]), .B(I_a[2]), .Z(n316) );
  GTECH_XNOR3 U327 ( .A(n325), .B(n327), .C(n322), .Z(n302) );
  GTECH_NOT U328 ( .A(n326), .Z(n322) );
  GTECH_OAI21 U329 ( .A(n343), .B(n344), .C(n345), .Z(n326) );
  GTECH_OAI21 U330 ( .A(n346), .B(n347), .C(n348), .Z(n345) );
  GTECH_NOT U331 ( .A(n349), .Z(n327) );
  GTECH_NAND2 U332 ( .A(I_b[3]), .B(I_a[3]), .Z(n349) );
  GTECH_NOT U333 ( .A(n323), .Z(n325) );
  GTECH_NAND2 U334 ( .A(I_b[2]), .B(I_a[4]), .Z(n323) );
  GTECH_ADD_ABC U335 ( .A(n350), .B(n351), .C(n352), .COUT(n300) );
  GTECH_NOT U336 ( .A(n353), .Z(n352) );
  GTECH_XNOR3 U337 ( .A(n354), .B(n355), .C(n356), .Z(n351) );
  GTECH_NOT U338 ( .A(n357), .Z(n301) );
  GTECH_XNOR3 U339 ( .A(n309), .B(n310), .C(n330), .Z(n357) );
  GTECH_NOT U340 ( .A(n311), .Z(n330) );
  GTECH_OAI21 U341 ( .A(n358), .B(n359), .C(n360), .Z(n311) );
  GTECH_OAI21 U342 ( .A(n354), .B(n356), .C(n355), .Z(n360) );
  GTECH_NOT U343 ( .A(n361), .Z(n310) );
  GTECH_NAND2 U344 ( .A(I_a[5]), .B(I_b[1]), .Z(n361) );
  GTECH_NOT U345 ( .A(n331), .Z(n309) );
  GTECH_NAND2 U346 ( .A(I_a[6]), .B(I_b[0]), .Z(n331) );
  GTECH_XNOR3 U347 ( .A(n362), .B(n306), .C(n363), .Z(N145) );
  GTECH_NOT U348 ( .A(n305), .Z(n363) );
  GTECH_XOR2 U349 ( .A(n364), .B(n342), .Z(n305) );
  GTECH_NOT U350 ( .A(n365), .Z(n342) );
  GTECH_NAND2 U351 ( .A(I_b[5]), .B(I_a[0]), .Z(n365) );
  GTECH_NAND2 U352 ( .A(I_b[4]), .B(I_a[1]), .Z(n364) );
  GTECH_NOT U353 ( .A(n337), .Z(n306) );
  GTECH_XOR2 U354 ( .A(n366), .B(n350), .Z(n337) );
  GTECH_ADD_ABC U355 ( .A(n367), .B(n368), .C(n369), .COUT(n350) );
  GTECH_XNOR3 U356 ( .A(n370), .B(n371), .C(n372), .Z(n368) );
  GTECH_OA22 U357 ( .A(n373), .B(n374), .C(n375), .D(n376), .Z(n367) );
  GTECH_AND2 U358 ( .A(n375), .B(n376), .Z(n373) );
  GTECH_XOR4 U359 ( .A(n355), .B(n358), .C(n353), .D(n354), .Z(n366) );
  GTECH_NOT U360 ( .A(n359), .Z(n354) );
  GTECH_NAND2 U361 ( .A(I_a[5]), .B(I_b[0]), .Z(n359) );
  GTECH_XNOR3 U362 ( .A(n346), .B(n348), .C(n343), .Z(n353) );
  GTECH_NOT U363 ( .A(n347), .Z(n343) );
  GTECH_OAI21 U364 ( .A(n377), .B(n378), .C(n379), .Z(n347) );
  GTECH_NOT U365 ( .A(n380), .Z(n348) );
  GTECH_NAND2 U366 ( .A(I_b[3]), .B(I_a[2]), .Z(n380) );
  GTECH_NOT U367 ( .A(n344), .Z(n346) );
  GTECH_NAND2 U368 ( .A(I_b[2]), .B(I_a[3]), .Z(n344) );
  GTECH_NOT U369 ( .A(n356), .Z(n358) );
  GTECH_OAI21 U370 ( .A(n381), .B(n382), .C(n383), .Z(n356) );
  GTECH_OAI21 U371 ( .A(n370), .B(n372), .C(n371), .Z(n383) );
  GTECH_NOT U372 ( .A(n382), .Z(n370) );
  GTECH_NOT U373 ( .A(n384), .Z(n355) );
  GTECH_NAND2 U374 ( .A(I_a[4]), .B(I_b[1]), .Z(n384) );
  GTECH_NOT U375 ( .A(n304), .Z(n362) );
  GTECH_NAND3 U376 ( .A(I_a[0]), .B(n385), .C(I_b[4]), .Z(n304) );
  GTECH_XOR2 U377 ( .A(n386), .B(n385), .Z(N144) );
  GTECH_XOR2 U378 ( .A(n387), .B(n388), .Z(n385) );
  GTECH_OA22 U379 ( .A(n375), .B(n376), .C(n389), .D(n374), .Z(n388) );
  GTECH_AND_NOT U380 ( .A(n375), .B(n390), .Z(n389) );
  GTECH_XOR4 U381 ( .A(n371), .B(n381), .C(n382), .D(n369), .Z(n387) );
  GTECH_XNOR3 U382 ( .A(n391), .B(n392), .C(n393), .Z(n369) );
  GTECH_NOT U383 ( .A(n379), .Z(n393) );
  GTECH_NAND3 U384 ( .A(I_b[2]), .B(I_a[1]), .C(n394), .Z(n379) );
  GTECH_NOT U385 ( .A(n378), .Z(n392) );
  GTECH_NAND2 U386 ( .A(I_b[3]), .B(I_a[1]), .Z(n378) );
  GTECH_NOT U387 ( .A(n377), .Z(n391) );
  GTECH_NAND2 U388 ( .A(I_b[2]), .B(I_a[2]), .Z(n377) );
  GTECH_NAND2 U389 ( .A(I_a[4]), .B(I_b[0]), .Z(n382) );
  GTECH_NOT U390 ( .A(n372), .Z(n381) );
  GTECH_OAI21 U391 ( .A(n395), .B(n396), .C(n397), .Z(n372) );
  GTECH_OAI21 U392 ( .A(n398), .B(n399), .C(n400), .Z(n397) );
  GTECH_NOT U393 ( .A(n401), .Z(n371) );
  GTECH_NAND2 U394 ( .A(I_a[3]), .B(I_b[1]), .Z(n401) );
  GTECH_AND2 U395 ( .A(I_b[4]), .B(I_a[0]), .Z(n386) );
  GTECH_XNOR3 U396 ( .A(n402), .B(n376), .C(n403), .Z(N143) );
  GTECH_NOT U397 ( .A(n375), .Z(n403) );
  GTECH_XOR2 U398 ( .A(n404), .B(n394), .Z(n375) );
  GTECH_NOT U399 ( .A(n405), .Z(n394) );
  GTECH_NAND2 U400 ( .A(I_b[3]), .B(I_a[0]), .Z(n405) );
  GTECH_NAND2 U401 ( .A(I_b[2]), .B(I_a[1]), .Z(n404) );
  GTECH_NOT U402 ( .A(n390), .Z(n376) );
  GTECH_XNOR3 U403 ( .A(n398), .B(n400), .C(n395), .Z(n390) );
  GTECH_NOT U404 ( .A(n399), .Z(n395) );
  GTECH_OAI21 U405 ( .A(n406), .B(n407), .C(n408), .Z(n399) );
  GTECH_NOT U406 ( .A(n409), .Z(n400) );
  GTECH_NAND2 U407 ( .A(I_b[1]), .B(I_a[2]), .Z(n409) );
  GTECH_NOT U408 ( .A(n396), .Z(n398) );
  GTECH_NAND2 U409 ( .A(I_b[0]), .B(I_a[3]), .Z(n396) );
  GTECH_NOT U410 ( .A(n374), .Z(n402) );
  GTECH_NAND3 U411 ( .A(I_a[0]), .B(n410), .C(I_b[2]), .Z(n374) );
  GTECH_XOR2 U412 ( .A(n411), .B(n410), .Z(N142) );
  GTECH_NOT U413 ( .A(n412), .Z(n410) );
  GTECH_XNOR3 U414 ( .A(n413), .B(n414), .C(n415), .Z(n412) );
  GTECH_NOT U415 ( .A(n408), .Z(n415) );
  GTECH_NAND3 U416 ( .A(n416), .B(I_b[0]), .C(I_a[1]), .Z(n408) );
  GTECH_NOT U417 ( .A(n406), .Z(n414) );
  GTECH_NAND2 U418 ( .A(I_a[1]), .B(I_b[1]), .Z(n406) );
  GTECH_NOT U419 ( .A(n407), .Z(n413) );
  GTECH_NAND2 U420 ( .A(I_b[0]), .B(I_a[2]), .Z(n407) );
  GTECH_AND2 U421 ( .A(I_b[2]), .B(I_a[0]), .Z(n411) );
  GTECH_XOR2 U422 ( .A(n416), .B(n417), .Z(N141) );
  GTECH_AND2 U423 ( .A(I_a[1]), .B(I_b[0]), .Z(n417) );
  GTECH_NOT U424 ( .A(n418), .Z(n416) );
  GTECH_NAND2 U425 ( .A(I_a[0]), .B(I_b[1]), .Z(n418) );
  GTECH_AND2 U426 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

