
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385;

  GTECH_MUX2 U143 ( .A(n282), .B(n283), .S(n284), .Z(sum[9]) );
  GTECH_ADD_AB U144 ( .A(n285), .B(n286), .S(n283) );
  GTECH_NOT U145 ( .A(n287), .Z(n285) );
  GTECH_XNOR2 U146 ( .A(n288), .B(n286), .Z(n282) );
  GTECH_AOI21 U147 ( .A(a[9]), .B(b[9]), .C(n289), .Z(n286) );
  GTECH_NAND2 U148 ( .A(n290), .B(n291), .Z(sum[8]) );
  GTECH_OAI21 U149 ( .A(n292), .B(n287), .C(n284), .Z(n290) );
  GTECH_MUX2 U150 ( .A(n293), .B(n294), .S(n295), .Z(sum[7]) );
  GTECH_XNOR2 U151 ( .A(n296), .B(n297), .Z(n294) );
  GTECH_AND2 U152 ( .A(n298), .B(n299), .Z(n296) );
  GTECH_AO21 U153 ( .A(n300), .B(n301), .C(n302), .Z(n299) );
  GTECH_ADD_AB U154 ( .A(n303), .B(n297), .S(n293) );
  GTECH_ADD_AB U155 ( .A(b[7]), .B(a[7]), .S(n297) );
  GTECH_OAI21 U156 ( .A(n304), .B(n298), .C(n305), .Z(sum[6]) );
  GTECH_MUX2 U157 ( .A(n306), .B(n307), .S(b[6]), .Z(n305) );
  GTECH_NAND2 U158 ( .A(n301), .B(n304), .Z(n307) );
  GTECH_XNOR2 U159 ( .A(n301), .B(n304), .Z(n306) );
  GTECH_OA21 U160 ( .A(n308), .B(n295), .C(n302), .Z(n304) );
  GTECH_OAI21 U161 ( .A(n309), .B(n310), .C(n311), .Z(n302) );
  GTECH_MUX2 U162 ( .A(n312), .B(n313), .S(n314), .Z(sum[5]) );
  GTECH_AND_NOT U163 ( .A(n311), .B(n309), .Z(n314) );
  GTECH_OAI21 U164 ( .A(a[4]), .B(n315), .C(n316), .Z(n313) );
  GTECH_AO21 U165 ( .A(n315), .B(a[4]), .C(b[4]), .Z(n316) );
  GTECH_AO21 U166 ( .A(n317), .B(n315), .C(n310), .Z(n312) );
  GTECH_ADD_AB U167 ( .A(n318), .B(n295), .S(sum[4]) );
  GTECH_MUX2 U168 ( .A(n319), .B(n320), .S(cin), .Z(sum[3]) );
  GTECH_ADD_AB U169 ( .A(n321), .B(n322), .S(n320) );
  GTECH_ADD_AB U170 ( .A(n323), .B(n322), .S(n319) );
  GTECH_ADD_AB U171 ( .A(b[3]), .B(a[3]), .S(n322) );
  GTECH_ADD_ABC U172 ( .A(a[2]), .B(n324), .C(b[2]), .COUT(n323) );
  GTECH_MUX2 U173 ( .A(n325), .B(n326), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U174 ( .A(n327), .B(n328), .Z(n326) );
  GTECH_XNOR2 U175 ( .A(n324), .B(n328), .Z(n325) );
  GTECH_XNOR2 U176 ( .A(b[2]), .B(a[2]), .Z(n328) );
  GTECH_OA21 U177 ( .A(n329), .B(n330), .C(n331), .Z(n324) );
  GTECH_MUX2 U178 ( .A(n332), .B(n333), .S(n334), .Z(sum[1]) );
  GTECH_AND_NOT U179 ( .A(n331), .B(n329), .Z(n334) );
  GTECH_OAI21 U180 ( .A(cin), .B(n330), .C(n335), .Z(n333) );
  GTECH_AO21 U181 ( .A(n335), .B(cin), .C(n330), .Z(n332) );
  GTECH_MUX2 U182 ( .A(n336), .B(n337), .S(n338), .Z(sum[15]) );
  GTECH_XNOR2 U183 ( .A(n339), .B(n340), .Z(n337) );
  GTECH_OA21 U184 ( .A(n341), .B(n342), .C(n343), .Z(n339) );
  GTECH_ADD_AB U185 ( .A(n344), .B(n340), .S(n336) );
  GTECH_ADD_AB U186 ( .A(b[15]), .B(a[15]), .S(n340) );
  GTECH_MUX2 U187 ( .A(n345), .B(n346), .S(n347), .Z(sum[14]) );
  GTECH_OA21 U188 ( .A(n348), .B(n338), .C(n342), .Z(n347) );
  GTECH_OA21 U189 ( .A(n349), .B(n350), .C(n351), .Z(n342) );
  GTECH_ADD_AB U190 ( .A(b[14]), .B(a[14]), .S(n346) );
  GTECH_OR_NOT U191 ( .A(n341), .B(n343), .Z(n345) );
  GTECH_MUX2 U192 ( .A(n352), .B(n353), .S(n354), .Z(sum[13]) );
  GTECH_OA21 U193 ( .A(n355), .B(n338), .C(n350), .Z(n354) );
  GTECH_ADD_AB U194 ( .A(b[13]), .B(a[13]), .S(n353) );
  GTECH_OR_NOT U195 ( .A(n349), .B(n351), .Z(n352) );
  GTECH_NAND2 U196 ( .A(n356), .B(n357), .Z(sum[12]) );
  GTECH_AO21 U197 ( .A(n350), .B(n358), .C(n338), .Z(n357) );
  GTECH_MUX2 U198 ( .A(n359), .B(n360), .S(n284), .Z(sum[11]) );
  GTECH_ADD_AB U199 ( .A(n361), .B(n362), .S(n360) );
  GTECH_XNOR2 U200 ( .A(n363), .B(n362), .Z(n359) );
  GTECH_ADD_AB U201 ( .A(b[11]), .B(a[11]), .S(n362) );
  GTECH_AND2 U202 ( .A(n364), .B(n365), .Z(n363) );
  GTECH_OAI21 U203 ( .A(b[10]), .B(a[10]), .C(n366), .Z(n365) );
  GTECH_OAI21 U204 ( .A(n367), .B(n364), .C(n368), .Z(sum[10]) );
  GTECH_MUX2 U205 ( .A(n369), .B(n370), .S(b[10]), .Z(n368) );
  GTECH_OR_NOT U206 ( .A(a[10]), .B(n367), .Z(n370) );
  GTECH_ADD_AB U207 ( .A(a[10]), .B(n367), .S(n369) );
  GTECH_AOI21 U208 ( .A(n371), .B(n284), .C(n366), .Z(n367) );
  GTECH_OAI2N2 U209 ( .A(n289), .B(n288), .C(a[9]), .D(b[9]), .Z(n366) );
  GTECH_NOT U210 ( .A(n292), .Z(n288) );
  GTECH_ADD_AB U211 ( .A(cin), .B(n372), .S(sum[0]) );
  GTECH_OAI21 U212 ( .A(n338), .B(n373), .C(n356), .Z(cout) );
  GTECH_NOT U213 ( .A(n374), .Z(n356) );
  GTECH_AND3 U214 ( .A(n358), .B(n350), .C(n338), .Z(n374) );
  GTECH_NAND2 U215 ( .A(b[12]), .B(a[12]), .Z(n350) );
  GTECH_AOI21 U216 ( .A(n344), .B(a[15]), .C(n375), .Z(n373) );
  GTECH_OA21 U217 ( .A(a[15]), .B(n344), .C(b[15]), .Z(n375) );
  GTECH_NAND2 U218 ( .A(n376), .B(n343), .Z(n344) );
  GTECH_NAND2 U219 ( .A(a[14]), .B(b[14]), .Z(n343) );
  GTECH_AO21 U220 ( .A(n348), .B(n351), .C(n341), .Z(n376) );
  GTECH_NOR2 U221 ( .A(b[14]), .B(a[14]), .Z(n341) );
  GTECH_NAND2 U222 ( .A(b[13]), .B(a[13]), .Z(n351) );
  GTECH_OR_NOT U223 ( .A(n349), .B(n358), .Z(n348) );
  GTECH_NOT U224 ( .A(n355), .Z(n358) );
  GTECH_NOR2 U225 ( .A(b[12]), .B(a[12]), .Z(n355) );
  GTECH_NOR2 U226 ( .A(a[13]), .B(b[13]), .Z(n349) );
  GTECH_OA21 U227 ( .A(n377), .B(n378), .C(n291), .Z(n338) );
  GTECH_OR3 U228 ( .A(n287), .B(n292), .C(n284), .Z(n291) );
  GTECH_NOT U229 ( .A(n378), .Z(n284) );
  GTECH_AND2 U230 ( .A(b[8]), .B(a[8]), .Z(n292) );
  GTECH_MUX2 U231 ( .A(n379), .B(n318), .S(n295), .Z(n378) );
  GTECH_NOT U232 ( .A(n315), .Z(n295) );
  GTECH_MUX2 U233 ( .A(n372), .B(n380), .S(cin), .Z(n315) );
  GTECH_OA21 U234 ( .A(a[3]), .B(n321), .C(n381), .Z(n380) );
  GTECH_AO21 U235 ( .A(n321), .B(a[3]), .C(b[3]), .Z(n381) );
  GTECH_ADD_ABC U236 ( .A(n327), .B(a[2]), .C(b[2]), .COUT(n321) );
  GTECH_OA21 U237 ( .A(n329), .B(n335), .C(n331), .Z(n327) );
  GTECH_OR2 U238 ( .A(b[1]), .B(a[1]), .Z(n331) );
  GTECH_AND2 U239 ( .A(b[1]), .B(a[1]), .Z(n329) );
  GTECH_AND_NOT U240 ( .A(n335), .B(n330), .Z(n372) );
  GTECH_AND2 U241 ( .A(b[0]), .B(a[0]), .Z(n330) );
  GTECH_OR2 U242 ( .A(b[0]), .B(a[0]), .Z(n335) );
  GTECH_OR_NOT U243 ( .A(n310), .B(n317), .Z(n318) );
  GTECH_AND2 U244 ( .A(a[4]), .B(b[4]), .Z(n310) );
  GTECH_AOI21 U245 ( .A(n303), .B(a[7]), .C(n382), .Z(n379) );
  GTECH_OA21 U246 ( .A(a[7]), .B(n303), .C(b[7]), .Z(n382) );
  GTECH_NAND2 U247 ( .A(n383), .B(n298), .Z(n303) );
  GTECH_OR_NOT U248 ( .A(n301), .B(b[6]), .Z(n298) );
  GTECH_AO21 U249 ( .A(n301), .B(n300), .C(n308), .Z(n383) );
  GTECH_OAI21 U250 ( .A(n309), .B(n317), .C(n311), .Z(n308) );
  GTECH_OR2 U251 ( .A(b[5]), .B(a[5]), .Z(n311) );
  GTECH_OR2 U252 ( .A(a[4]), .B(b[4]), .Z(n317) );
  GTECH_AND2 U253 ( .A(b[5]), .B(a[5]), .Z(n309) );
  GTECH_NOT U254 ( .A(b[6]), .Z(n300) );
  GTECH_NOT U255 ( .A(a[6]), .Z(n301) );
  GTECH_AOI21 U256 ( .A(n361), .B(a[11]), .C(n384), .Z(n377) );
  GTECH_OA21 U257 ( .A(a[11]), .B(n361), .C(b[11]), .Z(n384) );
  GTECH_NAND2 U258 ( .A(n385), .B(n364), .Z(n361) );
  GTECH_NAND2 U259 ( .A(a[10]), .B(b[10]), .Z(n364) );
  GTECH_OAI21 U260 ( .A(a[10]), .B(b[10]), .C(n371), .Z(n385) );
  GTECH_OAI2N2 U261 ( .A(n289), .B(n287), .C(a[9]), .D(b[9]), .Z(n371) );
  GTECH_NOR2 U262 ( .A(b[8]), .B(a[8]), .Z(n287) );
  GTECH_NOR2 U263 ( .A(b[9]), .B(a[9]), .Z(n289) );
endmodule

