
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI21 U82 ( .A(n93), .B(n94), .C(n95), .Z(n87) );
  GTECH_OAI21 U83 ( .A(n96), .B(n97), .C(n98), .Z(n95) );
  GTECH_NOT U84 ( .A(n93), .Z(n97) );
  GTECH_XOR2 U85 ( .A(n90), .B(n99), .Z(n86) );
  GTECH_NOT U86 ( .A(n89), .Z(n99) );
  GTECH_OAI21 U87 ( .A(n100), .B(n101), .C(n102), .Z(n89) );
  GTECH_OAI21 U88 ( .A(n103), .B(n104), .C(n105), .Z(n102) );
  GTECH_NAND2 U89 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n106), .Z(n84) );
  GTECH_NAND2 U91 ( .A(n107), .B(n108), .Z(n106) );
  GTECH_XOR2 U92 ( .A(n108), .B(n107), .Z(N153) );
  GTECH_NOT U93 ( .A(n109), .Z(n107) );
  GTECH_XNOR3 U94 ( .A(n96), .B(n93), .C(n110), .Z(n109) );
  GTECH_NOT U95 ( .A(n98), .Z(n110) );
  GTECH_XNOR3 U96 ( .A(n103), .B(n105), .C(n100), .Z(n98) );
  GTECH_NOT U97 ( .A(n104), .Z(n100) );
  GTECH_OAI21 U98 ( .A(n111), .B(n112), .C(n113), .Z(n104) );
  GTECH_OAI21 U99 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_NOT U100 ( .A(n117), .Z(n105) );
  GTECH_NAND2 U101 ( .A(I_b[7]), .B(I_a[6]), .Z(n117) );
  GTECH_NOT U102 ( .A(n101), .Z(n103) );
  GTECH_NAND2 U103 ( .A(I_a[7]), .B(I_b[6]), .Z(n101) );
  GTECH_ADD_ABC U104 ( .A(n118), .B(n119), .C(n120), .COUT(n93) );
  GTECH_NOT U105 ( .A(n121), .Z(n120) );
  GTECH_XOR2 U106 ( .A(n122), .B(n123), .Z(n119) );
  GTECH_AND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n123) );
  GTECH_NOT U108 ( .A(n94), .Z(n96) );
  GTECH_NAND2 U109 ( .A(I_a[7]), .B(n124), .Z(n94) );
  GTECH_NOT U110 ( .A(n125), .Z(n108) );
  GTECH_NAND2 U111 ( .A(n126), .B(n127), .Z(n125) );
  GTECH_NOT U112 ( .A(n128), .Z(n127) );
  GTECH_XOR2 U113 ( .A(n128), .B(n129), .Z(N152) );
  GTECH_NOT U114 ( .A(n126), .Z(n129) );
  GTECH_XOR4 U115 ( .A(n130), .B(n122), .C(n121), .D(n118), .Z(n126) );
  GTECH_ADD_ABC U116 ( .A(n131), .B(n132), .C(n133), .COUT(n118) );
  GTECH_XNOR3 U117 ( .A(n134), .B(n135), .C(n136), .Z(n132) );
  GTECH_XNOR3 U118 ( .A(n114), .B(n116), .C(n111), .Z(n121) );
  GTECH_NOT U119 ( .A(n115), .Z(n111) );
  GTECH_OAI21 U120 ( .A(n137), .B(n138), .C(n139), .Z(n115) );
  GTECH_OAI21 U121 ( .A(n140), .B(n141), .C(n142), .Z(n139) );
  GTECH_NOT U122 ( .A(n143), .Z(n116) );
  GTECH_NAND2 U123 ( .A(I_b[7]), .B(I_a[5]), .Z(n143) );
  GTECH_NOT U124 ( .A(n112), .Z(n114) );
  GTECH_NAND2 U125 ( .A(I_b[6]), .B(I_a[6]), .Z(n112) );
  GTECH_NOT U126 ( .A(n124), .Z(n122) );
  GTECH_OAI21 U127 ( .A(n144), .B(n145), .C(n146), .Z(n124) );
  GTECH_OAI21 U128 ( .A(n134), .B(n136), .C(n135), .Z(n146) );
  GTECH_AND2 U129 ( .A(I_a[7]), .B(I_b[5]), .Z(n130) );
  GTECH_ADD_ABC U130 ( .A(n147), .B(n148), .C(n149), .COUT(n128) );
  GTECH_OA22 U131 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n148) );
  GTECH_OA21 U132 ( .A(n154), .B(n155), .C(n156), .Z(n147) );
  GTECH_XNOR3 U133 ( .A(n157), .B(n149), .C(n158), .Z(N151) );
  GTECH_OA21 U134 ( .A(n154), .B(n155), .C(n156), .Z(n158) );
  GTECH_OAI21 U135 ( .A(n159), .B(n160), .C(n161), .Z(n156) );
  GTECH_XOR2 U136 ( .A(n131), .B(n162), .Z(n149) );
  GTECH_XOR4 U137 ( .A(n135), .B(n144), .C(n133), .D(n134), .Z(n162) );
  GTECH_NOT U138 ( .A(n145), .Z(n134) );
  GTECH_NAND2 U139 ( .A(I_a[7]), .B(I_b[4]), .Z(n145) );
  GTECH_NOT U140 ( .A(n163), .Z(n133) );
  GTECH_XNOR3 U141 ( .A(n140), .B(n142), .C(n137), .Z(n163) );
  GTECH_NOT U142 ( .A(n141), .Z(n137) );
  GTECH_OAI21 U143 ( .A(n164), .B(n165), .C(n166), .Z(n141) );
  GTECH_OAI21 U144 ( .A(n167), .B(n168), .C(n169), .Z(n166) );
  GTECH_NOT U145 ( .A(n170), .Z(n142) );
  GTECH_NAND2 U146 ( .A(I_b[7]), .B(I_a[4]), .Z(n170) );
  GTECH_NOT U147 ( .A(n138), .Z(n140) );
  GTECH_NAND2 U148 ( .A(I_b[6]), .B(I_a[5]), .Z(n138) );
  GTECH_NOT U149 ( .A(n136), .Z(n144) );
  GTECH_OAI21 U150 ( .A(n171), .B(n172), .C(n173), .Z(n136) );
  GTECH_OAI21 U151 ( .A(n174), .B(n175), .C(n176), .Z(n173) );
  GTECH_NOT U152 ( .A(n177), .Z(n135) );
  GTECH_NAND2 U153 ( .A(I_a[6]), .B(I_b[5]), .Z(n177) );
  GTECH_ADD_ABC U154 ( .A(n178), .B(n179), .C(n180), .COUT(n131) );
  GTECH_NOT U155 ( .A(n181), .Z(n180) );
  GTECH_XNOR3 U156 ( .A(n174), .B(n176), .C(n175), .Z(n179) );
  GTECH_OA22 U157 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n157) );
  GTECH_NOT U158 ( .A(n182), .Z(n153) );
  GTECH_NOT U159 ( .A(I_a[7]), .Z(n151) );
  GTECH_XNOR3 U160 ( .A(n154), .B(n159), .C(n161), .Z(N150) );
  GTECH_XOR2 U161 ( .A(n183), .B(n178), .Z(n161) );
  GTECH_ADD_ABC U162 ( .A(n184), .B(n185), .C(n186), .COUT(n178) );
  GTECH_NOT U163 ( .A(n187), .Z(n186) );
  GTECH_XNOR3 U164 ( .A(n188), .B(n189), .C(n190), .Z(n185) );
  GTECH_XOR4 U165 ( .A(n176), .B(n171), .C(n181), .D(n174), .Z(n183) );
  GTECH_NOT U166 ( .A(n172), .Z(n174) );
  GTECH_NAND2 U167 ( .A(I_a[6]), .B(I_b[4]), .Z(n172) );
  GTECH_XNOR3 U168 ( .A(n167), .B(n169), .C(n164), .Z(n181) );
  GTECH_NOT U169 ( .A(n168), .Z(n164) );
  GTECH_OAI21 U170 ( .A(n191), .B(n192), .C(n193), .Z(n168) );
  GTECH_OAI21 U171 ( .A(n194), .B(n195), .C(n196), .Z(n193) );
  GTECH_NOT U172 ( .A(n197), .Z(n169) );
  GTECH_NAND2 U173 ( .A(I_b[7]), .B(I_a[3]), .Z(n197) );
  GTECH_NOT U174 ( .A(n165), .Z(n167) );
  GTECH_NAND2 U175 ( .A(I_b[6]), .B(I_a[4]), .Z(n165) );
  GTECH_NOT U176 ( .A(n175), .Z(n171) );
  GTECH_OAI21 U177 ( .A(n198), .B(n199), .C(n200), .Z(n175) );
  GTECH_OAI21 U178 ( .A(n188), .B(n190), .C(n189), .Z(n200) );
  GTECH_NOT U179 ( .A(n201), .Z(n176) );
  GTECH_NAND2 U180 ( .A(I_a[5]), .B(I_b[5]), .Z(n201) );
  GTECH_NOT U181 ( .A(n155), .Z(n159) );
  GTECH_XOR2 U182 ( .A(n182), .B(n152), .Z(n155) );
  GTECH_AOI2N2 U183 ( .A(n202), .B(n203), .C(n204), .D(n205), .Z(n152) );
  GTECH_NAND2 U184 ( .A(n204), .B(n205), .Z(n203) );
  GTECH_XOR2 U185 ( .A(n206), .B(n150), .Z(n182) );
  GTECH_OA21 U186 ( .A(n207), .B(n208), .C(n209), .Z(n150) );
  GTECH_OAI21 U187 ( .A(n210), .B(n211), .C(n212), .Z(n209) );
  GTECH_NAND2 U188 ( .A(I_a[7]), .B(I_b[3]), .Z(n206) );
  GTECH_NOT U189 ( .A(n160), .Z(n154) );
  GTECH_OAI21 U190 ( .A(n213), .B(n214), .C(n215), .Z(n160) );
  GTECH_OAI21 U191 ( .A(n216), .B(n217), .C(n218), .Z(n215) );
  GTECH_NOT U192 ( .A(n213), .Z(n217) );
  GTECH_XNOR3 U193 ( .A(n213), .B(n216), .C(n218), .Z(N149) );
  GTECH_XOR2 U194 ( .A(n219), .B(n184), .Z(n218) );
  GTECH_ADD_ABC U195 ( .A(n220), .B(n221), .C(n222), .COUT(n184) );
  GTECH_XNOR3 U196 ( .A(n223), .B(n224), .C(n225), .Z(n221) );
  GTECH_OA21 U197 ( .A(n226), .B(n227), .C(n228), .Z(n220) );
  GTECH_XOR4 U198 ( .A(n189), .B(n198), .C(n187), .D(n188), .Z(n219) );
  GTECH_NOT U199 ( .A(n199), .Z(n188) );
  GTECH_NAND2 U200 ( .A(I_a[5]), .B(I_b[4]), .Z(n199) );
  GTECH_XNOR3 U201 ( .A(n194), .B(n196), .C(n191), .Z(n187) );
  GTECH_NOT U202 ( .A(n195), .Z(n191) );
  GTECH_OAI21 U203 ( .A(n229), .B(n230), .C(n231), .Z(n195) );
  GTECH_NOT U204 ( .A(n232), .Z(n196) );
  GTECH_NAND2 U205 ( .A(I_b[7]), .B(I_a[2]), .Z(n232) );
  GTECH_NOT U206 ( .A(n192), .Z(n194) );
  GTECH_NAND2 U207 ( .A(I_b[6]), .B(I_a[3]), .Z(n192) );
  GTECH_NOT U208 ( .A(n190), .Z(n198) );
  GTECH_OAI21 U209 ( .A(n233), .B(n234), .C(n235), .Z(n190) );
  GTECH_OAI21 U210 ( .A(n223), .B(n225), .C(n224), .Z(n235) );
  GTECH_NOT U211 ( .A(n236), .Z(n189) );
  GTECH_NAND2 U212 ( .A(I_b[5]), .B(I_a[4]), .Z(n236) );
  GTECH_NOT U213 ( .A(n214), .Z(n216) );
  GTECH_XNOR3 U214 ( .A(n237), .B(n204), .C(n238), .Z(n214) );
  GTECH_NOT U215 ( .A(n202), .Z(n238) );
  GTECH_XNOR3 U216 ( .A(n210), .B(n212), .C(n207), .Z(n202) );
  GTECH_NOT U217 ( .A(n211), .Z(n207) );
  GTECH_OAI21 U218 ( .A(n239), .B(n240), .C(n241), .Z(n211) );
  GTECH_OAI21 U219 ( .A(n242), .B(n243), .C(n244), .Z(n241) );
  GTECH_NOT U220 ( .A(n245), .Z(n212) );
  GTECH_NAND2 U221 ( .A(I_a[6]), .B(I_b[3]), .Z(n245) );
  GTECH_NOT U222 ( .A(n208), .Z(n210) );
  GTECH_NAND2 U223 ( .A(I_a[7]), .B(I_b[2]), .Z(n208) );
  GTECH_ADD_ABC U224 ( .A(n246), .B(n247), .C(n248), .COUT(n204) );
  GTECH_NOT U225 ( .A(n249), .Z(n248) );
  GTECH_XOR2 U226 ( .A(n250), .B(n251), .Z(n247) );
  GTECH_AND2 U227 ( .A(I_a[7]), .B(I_b[1]), .Z(n251) );
  GTECH_NOT U228 ( .A(n205), .Z(n237) );
  GTECH_NAND2 U229 ( .A(I_a[7]), .B(n252), .Z(n205) );
  GTECH_ADD_ABC U230 ( .A(n253), .B(n254), .C(n255), .COUT(n213) );
  GTECH_XNOR3 U231 ( .A(n246), .B(n256), .C(n249), .Z(n254) );
  GTECH_XOR2 U232 ( .A(n257), .B(n253), .Z(N148) );
  GTECH_ADD_ABC U233 ( .A(n258), .B(n259), .C(n260), .COUT(n253) );
  GTECH_NOT U234 ( .A(n261), .Z(n260) );
  GTECH_XNOR3 U235 ( .A(n262), .B(n263), .C(n264), .Z(n259) );
  GTECH_XOR4 U236 ( .A(n256), .B(n246), .C(n249), .D(n255), .Z(n257) );
  GTECH_XOR2 U237 ( .A(n265), .B(n266), .Z(n255) );
  GTECH_XOR4 U238 ( .A(n224), .B(n233), .C(n222), .D(n223), .Z(n266) );
  GTECH_NOT U239 ( .A(n234), .Z(n223) );
  GTECH_NAND2 U240 ( .A(I_b[4]), .B(I_a[4]), .Z(n234) );
  GTECH_XNOR3 U241 ( .A(n267), .B(n268), .C(n269), .Z(n222) );
  GTECH_NOT U242 ( .A(n231), .Z(n269) );
  GTECH_NAND3 U243 ( .A(I_b[6]), .B(I_a[1]), .C(n270), .Z(n231) );
  GTECH_NOT U244 ( .A(n230), .Z(n268) );
  GTECH_NAND2 U245 ( .A(I_b[7]), .B(I_a[1]), .Z(n230) );
  GTECH_NOT U246 ( .A(n229), .Z(n267) );
  GTECH_NAND2 U247 ( .A(I_b[6]), .B(I_a[2]), .Z(n229) );
  GTECH_NOT U248 ( .A(n225), .Z(n233) );
  GTECH_OAI21 U249 ( .A(n271), .B(n272), .C(n273), .Z(n225) );
  GTECH_OAI21 U250 ( .A(n274), .B(n275), .C(n276), .Z(n273) );
  GTECH_NOT U251 ( .A(n277), .Z(n224) );
  GTECH_NAND2 U252 ( .A(I_b[5]), .B(I_a[3]), .Z(n277) );
  GTECH_OA21 U253 ( .A(n226), .B(n227), .C(n228), .Z(n265) );
  GTECH_OAI21 U254 ( .A(n278), .B(n279), .C(n280), .Z(n228) );
  GTECH_XNOR3 U255 ( .A(n242), .B(n244), .C(n239), .Z(n249) );
  GTECH_NOT U256 ( .A(n243), .Z(n239) );
  GTECH_OAI21 U257 ( .A(n281), .B(n282), .C(n283), .Z(n243) );
  GTECH_OAI21 U258 ( .A(n284), .B(n285), .C(n286), .Z(n283) );
  GTECH_NOT U259 ( .A(n287), .Z(n244) );
  GTECH_NAND2 U260 ( .A(I_a[5]), .B(I_b[3]), .Z(n287) );
  GTECH_NOT U261 ( .A(n240), .Z(n242) );
  GTECH_NAND2 U262 ( .A(I_a[6]), .B(I_b[2]), .Z(n240) );
  GTECH_ADD_ABC U263 ( .A(n262), .B(n288), .C(n289), .COUT(n246) );
  GTECH_XNOR3 U264 ( .A(n290), .B(n291), .C(n292), .Z(n288) );
  GTECH_XOR2 U265 ( .A(n293), .B(n250), .Z(n256) );
  GTECH_NOT U266 ( .A(n252), .Z(n250) );
  GTECH_OAI21 U267 ( .A(n294), .B(n295), .C(n296), .Z(n252) );
  GTECH_OAI21 U268 ( .A(n290), .B(n292), .C(n291), .Z(n296) );
  GTECH_AND2 U269 ( .A(I_a[7]), .B(I_b[1]), .Z(n293) );
  GTECH_XOR2 U270 ( .A(n297), .B(n258), .Z(N147) );
  GTECH_ADD_ABC U271 ( .A(n298), .B(n299), .C(n300), .COUT(n258) );
  GTECH_XNOR3 U272 ( .A(n301), .B(n302), .C(n303), .Z(n299) );
  GTECH_OA21 U273 ( .A(n304), .B(n305), .C(n306), .Z(n298) );
  GTECH_XOR4 U274 ( .A(n263), .B(n289), .C(n261), .D(n262), .Z(n297) );
  GTECH_ADD_ABC U275 ( .A(n301), .B(n307), .C(n308), .COUT(n262) );
  GTECH_NOT U276 ( .A(n303), .Z(n308) );
  GTECH_XNOR3 U277 ( .A(n309), .B(n310), .C(n311), .Z(n307) );
  GTECH_XNOR3 U278 ( .A(n280), .B(n227), .C(n279), .Z(n261) );
  GTECH_NOT U279 ( .A(n226), .Z(n279) );
  GTECH_XOR2 U280 ( .A(n312), .B(n270), .Z(n226) );
  GTECH_NOT U281 ( .A(n313), .Z(n270) );
  GTECH_NAND2 U282 ( .A(I_b[7]), .B(I_a[0]), .Z(n313) );
  GTECH_NAND2 U283 ( .A(I_b[6]), .B(I_a[1]), .Z(n312) );
  GTECH_NOT U284 ( .A(n278), .Z(n227) );
  GTECH_XNOR3 U285 ( .A(n274), .B(n276), .C(n271), .Z(n278) );
  GTECH_NOT U286 ( .A(n275), .Z(n271) );
  GTECH_OAI21 U287 ( .A(n314), .B(n315), .C(n316), .Z(n275) );
  GTECH_NOT U288 ( .A(n317), .Z(n276) );
  GTECH_NAND2 U289 ( .A(I_b[5]), .B(I_a[2]), .Z(n317) );
  GTECH_NOT U290 ( .A(n272), .Z(n274) );
  GTECH_NAND2 U291 ( .A(I_b[4]), .B(I_a[3]), .Z(n272) );
  GTECH_NOT U292 ( .A(n318), .Z(n280) );
  GTECH_NAND3 U293 ( .A(I_a[0]), .B(n319), .C(I_b[6]), .Z(n318) );
  GTECH_NOT U294 ( .A(n320), .Z(n319) );
  GTECH_NOT U295 ( .A(n264), .Z(n289) );
  GTECH_XNOR3 U296 ( .A(n284), .B(n286), .C(n281), .Z(n264) );
  GTECH_NOT U297 ( .A(n285), .Z(n281) );
  GTECH_OAI21 U298 ( .A(n321), .B(n322), .C(n323), .Z(n285) );
  GTECH_OAI21 U299 ( .A(n324), .B(n325), .C(n326), .Z(n323) );
  GTECH_NOT U300 ( .A(n327), .Z(n286) );
  GTECH_NAND2 U301 ( .A(I_b[3]), .B(I_a[4]), .Z(n327) );
  GTECH_NOT U302 ( .A(n282), .Z(n284) );
  GTECH_NAND2 U303 ( .A(I_a[5]), .B(I_b[2]), .Z(n282) );
  GTECH_NOT U304 ( .A(n328), .Z(n263) );
  GTECH_XNOR3 U305 ( .A(n290), .B(n291), .C(n294), .Z(n328) );
  GTECH_NOT U306 ( .A(n292), .Z(n294) );
  GTECH_OAI21 U307 ( .A(n329), .B(n330), .C(n331), .Z(n292) );
  GTECH_OAI21 U308 ( .A(n309), .B(n311), .C(n310), .Z(n331) );
  GTECH_NOT U309 ( .A(n332), .Z(n291) );
  GTECH_NAND2 U310 ( .A(I_a[6]), .B(I_b[1]), .Z(n332) );
  GTECH_NOT U311 ( .A(n295), .Z(n290) );
  GTECH_NAND2 U312 ( .A(I_a[7]), .B(I_b[0]), .Z(n295) );
  GTECH_XOR2 U313 ( .A(n333), .B(n334), .Z(N146) );
  GTECH_OA21 U314 ( .A(n304), .B(n305), .C(n306), .Z(n334) );
  GTECH_OAI21 U315 ( .A(n335), .B(n336), .C(n337), .Z(n306) );
  GTECH_XOR4 U316 ( .A(n302), .B(n301), .C(n303), .D(n300), .Z(n333) );
  GTECH_XOR2 U317 ( .A(n320), .B(n338), .Z(n300) );
  GTECH_AND2 U318 ( .A(I_b[6]), .B(I_a[0]), .Z(n338) );
  GTECH_XNOR3 U319 ( .A(n339), .B(n340), .C(n341), .Z(n320) );
  GTECH_NOT U320 ( .A(n316), .Z(n341) );
  GTECH_NAND3 U321 ( .A(I_b[4]), .B(I_a[1]), .C(n342), .Z(n316) );
  GTECH_NOT U322 ( .A(n315), .Z(n340) );
  GTECH_NAND2 U323 ( .A(I_b[5]), .B(I_a[1]), .Z(n315) );
  GTECH_NOT U324 ( .A(n314), .Z(n339) );
  GTECH_NAND2 U325 ( .A(I_b[4]), .B(I_a[2]), .Z(n314) );
  GTECH_XNOR3 U326 ( .A(n324), .B(n326), .C(n321), .Z(n303) );
  GTECH_NOT U327 ( .A(n325), .Z(n321) );
  GTECH_OAI21 U328 ( .A(n343), .B(n344), .C(n345), .Z(n325) );
  GTECH_OAI21 U329 ( .A(n346), .B(n347), .C(n348), .Z(n345) );
  GTECH_NOT U330 ( .A(n349), .Z(n326) );
  GTECH_NAND2 U331 ( .A(I_b[3]), .B(I_a[3]), .Z(n349) );
  GTECH_NOT U332 ( .A(n322), .Z(n324) );
  GTECH_NAND2 U333 ( .A(I_b[2]), .B(I_a[4]), .Z(n322) );
  GTECH_ADD_ABC U334 ( .A(n350), .B(n351), .C(n352), .COUT(n301) );
  GTECH_NOT U335 ( .A(n353), .Z(n352) );
  GTECH_XNOR3 U336 ( .A(n354), .B(n355), .C(n356), .Z(n351) );
  GTECH_NOT U337 ( .A(n357), .Z(n302) );
  GTECH_XNOR3 U338 ( .A(n309), .B(n310), .C(n329), .Z(n357) );
  GTECH_NOT U339 ( .A(n311), .Z(n329) );
  GTECH_OAI21 U340 ( .A(n358), .B(n359), .C(n360), .Z(n311) );
  GTECH_OAI21 U341 ( .A(n354), .B(n356), .C(n355), .Z(n360) );
  GTECH_NOT U342 ( .A(n361), .Z(n310) );
  GTECH_NAND2 U343 ( .A(I_a[5]), .B(I_b[1]), .Z(n361) );
  GTECH_NOT U344 ( .A(n330), .Z(n309) );
  GTECH_NAND2 U345 ( .A(I_a[6]), .B(I_b[0]), .Z(n330) );
  GTECH_XNOR3 U346 ( .A(n337), .B(n305), .C(n336), .Z(N145) );
  GTECH_NOT U347 ( .A(n304), .Z(n336) );
  GTECH_XOR2 U348 ( .A(n362), .B(n342), .Z(n304) );
  GTECH_NOT U349 ( .A(n363), .Z(n342) );
  GTECH_NAND2 U350 ( .A(I_b[5]), .B(I_a[0]), .Z(n363) );
  GTECH_NAND2 U351 ( .A(I_b[4]), .B(I_a[1]), .Z(n362) );
  GTECH_NOT U352 ( .A(n335), .Z(n305) );
  GTECH_XOR2 U353 ( .A(n364), .B(n350), .Z(n335) );
  GTECH_ADD_ABC U354 ( .A(n365), .B(n366), .C(n367), .COUT(n350) );
  GTECH_XNOR3 U355 ( .A(n368), .B(n369), .C(n370), .Z(n366) );
  GTECH_OA21 U356 ( .A(n371), .B(n372), .C(n373), .Z(n365) );
  GTECH_XOR4 U357 ( .A(n355), .B(n358), .C(n353), .D(n354), .Z(n364) );
  GTECH_NOT U358 ( .A(n359), .Z(n354) );
  GTECH_NAND2 U359 ( .A(I_a[5]), .B(I_b[0]), .Z(n359) );
  GTECH_XNOR3 U360 ( .A(n346), .B(n348), .C(n343), .Z(n353) );
  GTECH_NOT U361 ( .A(n347), .Z(n343) );
  GTECH_OAI21 U362 ( .A(n374), .B(n375), .C(n376), .Z(n347) );
  GTECH_NOT U363 ( .A(n377), .Z(n348) );
  GTECH_NAND2 U364 ( .A(I_b[3]), .B(I_a[2]), .Z(n377) );
  GTECH_NOT U365 ( .A(n344), .Z(n346) );
  GTECH_NAND2 U366 ( .A(I_b[2]), .B(I_a[3]), .Z(n344) );
  GTECH_NOT U367 ( .A(n356), .Z(n358) );
  GTECH_OAI21 U368 ( .A(n378), .B(n379), .C(n380), .Z(n356) );
  GTECH_OAI21 U369 ( .A(n368), .B(n370), .C(n369), .Z(n380) );
  GTECH_NOT U370 ( .A(n379), .Z(n368) );
  GTECH_NOT U371 ( .A(n381), .Z(n355) );
  GTECH_NAND2 U372 ( .A(I_a[4]), .B(I_b[1]), .Z(n381) );
  GTECH_NOT U373 ( .A(n382), .Z(n337) );
  GTECH_NAND3 U374 ( .A(I_a[0]), .B(n383), .C(I_b[4]), .Z(n382) );
  GTECH_XOR2 U375 ( .A(n384), .B(n383), .Z(N144) );
  GTECH_XOR2 U376 ( .A(n385), .B(n386), .Z(n383) );
  GTECH_OA21 U377 ( .A(n371), .B(n372), .C(n373), .Z(n386) );
  GTECH_OAI21 U378 ( .A(n387), .B(n388), .C(n389), .Z(n373) );
  GTECH_XOR4 U379 ( .A(n369), .B(n378), .C(n379), .D(n367), .Z(n385) );
  GTECH_XNOR3 U380 ( .A(n390), .B(n391), .C(n392), .Z(n367) );
  GTECH_NOT U381 ( .A(n376), .Z(n392) );
  GTECH_NAND3 U382 ( .A(I_b[2]), .B(I_a[1]), .C(n393), .Z(n376) );
  GTECH_NOT U383 ( .A(n375), .Z(n391) );
  GTECH_NAND2 U384 ( .A(I_b[3]), .B(I_a[1]), .Z(n375) );
  GTECH_NOT U385 ( .A(n374), .Z(n390) );
  GTECH_NAND2 U386 ( .A(I_b[2]), .B(I_a[2]), .Z(n374) );
  GTECH_NAND2 U387 ( .A(I_a[4]), .B(I_b[0]), .Z(n379) );
  GTECH_NOT U388 ( .A(n370), .Z(n378) );
  GTECH_OAI21 U389 ( .A(n394), .B(n395), .C(n396), .Z(n370) );
  GTECH_OAI21 U390 ( .A(n397), .B(n398), .C(n399), .Z(n396) );
  GTECH_NOT U391 ( .A(n400), .Z(n369) );
  GTECH_NAND2 U392 ( .A(I_a[3]), .B(I_b[1]), .Z(n400) );
  GTECH_AND2 U393 ( .A(I_b[4]), .B(I_a[0]), .Z(n384) );
  GTECH_XNOR3 U394 ( .A(n389), .B(n372), .C(n388), .Z(N143) );
  GTECH_NOT U395 ( .A(n371), .Z(n388) );
  GTECH_XOR2 U396 ( .A(n401), .B(n393), .Z(n371) );
  GTECH_NOT U397 ( .A(n402), .Z(n393) );
  GTECH_NAND2 U398 ( .A(I_b[3]), .B(I_a[0]), .Z(n402) );
  GTECH_NAND2 U399 ( .A(I_b[2]), .B(I_a[1]), .Z(n401) );
  GTECH_NOT U400 ( .A(n387), .Z(n372) );
  GTECH_XNOR3 U401 ( .A(n397), .B(n399), .C(n394), .Z(n387) );
  GTECH_NOT U402 ( .A(n398), .Z(n394) );
  GTECH_OAI21 U403 ( .A(n403), .B(n404), .C(n405), .Z(n398) );
  GTECH_NOT U404 ( .A(n406), .Z(n399) );
  GTECH_NAND2 U405 ( .A(I_b[1]), .B(I_a[2]), .Z(n406) );
  GTECH_NOT U406 ( .A(n395), .Z(n397) );
  GTECH_NAND2 U407 ( .A(I_b[0]), .B(I_a[3]), .Z(n395) );
  GTECH_NOT U408 ( .A(n407), .Z(n389) );
  GTECH_NAND3 U409 ( .A(I_a[0]), .B(n408), .C(I_b[2]), .Z(n407) );
  GTECH_XOR2 U410 ( .A(n409), .B(n408), .Z(N142) );
  GTECH_NOT U411 ( .A(n410), .Z(n408) );
  GTECH_XNOR3 U412 ( .A(n411), .B(n412), .C(n413), .Z(n410) );
  GTECH_NOT U413 ( .A(n405), .Z(n413) );
  GTECH_NAND3 U414 ( .A(n414), .B(I_b[0]), .C(I_a[1]), .Z(n405) );
  GTECH_NOT U415 ( .A(n403), .Z(n412) );
  GTECH_NAND2 U416 ( .A(I_a[1]), .B(I_b[1]), .Z(n403) );
  GTECH_NOT U417 ( .A(n404), .Z(n411) );
  GTECH_NAND2 U418 ( .A(I_b[0]), .B(I_a[2]), .Z(n404) );
  GTECH_AND2 U419 ( .A(I_b[2]), .B(I_a[0]), .Z(n409) );
  GTECH_XOR2 U420 ( .A(n414), .B(n415), .Z(N141) );
  GTECH_AND2 U421 ( .A(I_a[1]), .B(I_b[0]), .Z(n415) );
  GTECH_NOT U422 ( .A(n416), .Z(n414) );
  GTECH_NAND2 U423 ( .A(I_a[0]), .B(I_b[1]), .Z(n416) );
  GTECH_AND2 U424 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

