
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_OAI21 U75 ( .A(n83), .B(n84), .C(n85), .Z(N155) );
  GTECH_OA22 U76 ( .A(n86), .B(n87), .C(n88), .D(n89), .Z(n85) );
  GTECH_NOT U77 ( .A(n90), .Z(n87) );
  GTECH_XOR2 U78 ( .A(n91), .B(n92), .Z(N154) );
  GTECH_NOT U79 ( .A(n83), .Z(n92) );
  GTECH_XOR2 U80 ( .A(n90), .B(n86), .Z(n83) );
  GTECH_AOI2N2 U81 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n86) );
  GTECH_NAND2 U82 ( .A(n95), .B(n96), .Z(n94) );
  GTECH_XOR2 U83 ( .A(n89), .B(n88), .Z(n90) );
  GTECH_AND2 U84 ( .A(n97), .B(n98), .Z(n88) );
  GTECH_OR_NOT U85 ( .A(n99), .B(n100), .Z(n98) );
  GTECH_OAI21 U86 ( .A(n101), .B(n100), .C(n102), .Z(n97) );
  GTECH_NAND2 U87 ( .A(I_b[7]), .B(I_a[7]), .Z(n89) );
  GTECH_NOT U88 ( .A(n84), .Z(n91) );
  GTECH_NAND2 U89 ( .A(n103), .B(n104), .Z(n84) );
  GTECH_XOR2 U90 ( .A(n104), .B(n103), .Z(N153) );
  GTECH_NOT U91 ( .A(n105), .Z(n103) );
  GTECH_XOR3 U92 ( .A(n106), .B(n95), .C(n93), .Z(n105) );
  GTECH_XOR3 U93 ( .A(n101), .B(n102), .C(n100), .Z(n93) );
  GTECH_OAI21 U94 ( .A(n107), .B(n108), .C(n109), .Z(n100) );
  GTECH_OAI21 U95 ( .A(n110), .B(n111), .C(n112), .Z(n109) );
  GTECH_NOT U96 ( .A(n111), .Z(n107) );
  GTECH_NOT U97 ( .A(n113), .Z(n102) );
  GTECH_NAND2 U98 ( .A(I_b[7]), .B(I_a[6]), .Z(n113) );
  GTECH_NOT U99 ( .A(n99), .Z(n101) );
  GTECH_NAND2 U100 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U101 ( .A(n114), .B(n115), .C(n116), .COUT(n95) );
  GTECH_NOT U102 ( .A(n117), .Z(n116) );
  GTECH_XOR2 U103 ( .A(n118), .B(n119), .Z(n115) );
  GTECH_AND2 U104 ( .A(I_a[7]), .B(I_b[5]), .Z(n119) );
  GTECH_NOT U105 ( .A(n120), .Z(n118) );
  GTECH_NOT U106 ( .A(n96), .Z(n106) );
  GTECH_NAND2 U107 ( .A(I_a[7]), .B(n120), .Z(n96) );
  GTECH_NOT U108 ( .A(n121), .Z(n104) );
  GTECH_NAND2 U109 ( .A(n122), .B(n123), .Z(n121) );
  GTECH_NOT U110 ( .A(n124), .Z(n123) );
  GTECH_XOR2 U111 ( .A(n124), .B(n125), .Z(N152) );
  GTECH_NOT U112 ( .A(n122), .Z(n125) );
  GTECH_XNOR4 U113 ( .A(n126), .B(n117), .C(n120), .D(n114), .Z(n122) );
  GTECH_ADD_ABC U114 ( .A(n127), .B(n128), .C(n129), .COUT(n114) );
  GTECH_NOT U115 ( .A(n130), .Z(n129) );
  GTECH_XOR3 U116 ( .A(n131), .B(n132), .C(n133), .Z(n128) );
  GTECH_OAI21 U117 ( .A(n133), .B(n134), .C(n135), .Z(n120) );
  GTECH_OAI21 U118 ( .A(n131), .B(n136), .C(n132), .Z(n135) );
  GTECH_NOT U119 ( .A(n136), .Z(n133) );
  GTECH_XOR3 U120 ( .A(n110), .B(n112), .C(n111), .Z(n117) );
  GTECH_OAI21 U121 ( .A(n137), .B(n138), .C(n139), .Z(n111) );
  GTECH_OAI21 U122 ( .A(n140), .B(n141), .C(n142), .Z(n139) );
  GTECH_NOT U123 ( .A(n141), .Z(n137) );
  GTECH_NOT U124 ( .A(n143), .Z(n112) );
  GTECH_NAND2 U125 ( .A(I_b[7]), .B(I_a[5]), .Z(n143) );
  GTECH_NOT U126 ( .A(n108), .Z(n110) );
  GTECH_NAND2 U127 ( .A(I_b[6]), .B(I_a[6]), .Z(n108) );
  GTECH_AND2 U128 ( .A(I_a[7]), .B(I_b[5]), .Z(n126) );
  GTECH_ADD_ABC U129 ( .A(n144), .B(n145), .C(n146), .COUT(n124) );
  GTECH_NOT U130 ( .A(n147), .Z(n146) );
  GTECH_OA22 U131 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n145) );
  GTECH_OA21 U132 ( .A(n152), .B(n153), .C(n154), .Z(n144) );
  GTECH_XOR3 U133 ( .A(n155), .B(n147), .C(n156), .Z(N151) );
  GTECH_OA21 U134 ( .A(n152), .B(n153), .C(n154), .Z(n156) );
  GTECH_OAI21 U135 ( .A(n157), .B(n158), .C(n159), .Z(n154) );
  GTECH_XOR2 U136 ( .A(n160), .B(n127), .Z(n147) );
  GTECH_ADD_ABC U137 ( .A(n161), .B(n162), .C(n163), .COUT(n127) );
  GTECH_NOT U138 ( .A(n164), .Z(n163) );
  GTECH_XOR3 U139 ( .A(n165), .B(n166), .C(n167), .Z(n162) );
  GTECH_XNOR4 U140 ( .A(n132), .B(n136), .C(n130), .D(n131), .Z(n160) );
  GTECH_NOT U141 ( .A(n134), .Z(n131) );
  GTECH_NAND2 U142 ( .A(I_a[7]), .B(I_b[4]), .Z(n134) );
  GTECH_XOR3 U143 ( .A(n140), .B(n142), .C(n141), .Z(n130) );
  GTECH_OAI21 U144 ( .A(n168), .B(n169), .C(n170), .Z(n141) );
  GTECH_OAI21 U145 ( .A(n171), .B(n172), .C(n173), .Z(n170) );
  GTECH_NOT U146 ( .A(n172), .Z(n168) );
  GTECH_NOT U147 ( .A(n174), .Z(n142) );
  GTECH_NAND2 U148 ( .A(I_b[7]), .B(I_a[4]), .Z(n174) );
  GTECH_NOT U149 ( .A(n138), .Z(n140) );
  GTECH_NAND2 U150 ( .A(I_b[6]), .B(I_a[5]), .Z(n138) );
  GTECH_OAI21 U151 ( .A(n167), .B(n175), .C(n176), .Z(n136) );
  GTECH_OAI21 U152 ( .A(n165), .B(n177), .C(n166), .Z(n176) );
  GTECH_NOT U153 ( .A(n177), .Z(n167) );
  GTECH_NOT U154 ( .A(n178), .Z(n132) );
  GTECH_NAND2 U155 ( .A(I_a[6]), .B(I_b[5]), .Z(n178) );
  GTECH_OA22 U156 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n155) );
  GTECH_NOT U157 ( .A(n179), .Z(n151) );
  GTECH_NOT U158 ( .A(I_a[7]), .Z(n149) );
  GTECH_XOR3 U159 ( .A(n152), .B(n157), .C(n180), .Z(N150) );
  GTECH_NOT U160 ( .A(n159), .Z(n180) );
  GTECH_XOR2 U161 ( .A(n181), .B(n161), .Z(n159) );
  GTECH_ADD_ABC U162 ( .A(n182), .B(n183), .C(n184), .COUT(n161) );
  GTECH_NOT U163 ( .A(n185), .Z(n184) );
  GTECH_XOR3 U164 ( .A(n186), .B(n187), .C(n188), .Z(n183) );
  GTECH_XNOR4 U165 ( .A(n166), .B(n177), .C(n164), .D(n165), .Z(n181) );
  GTECH_NOT U166 ( .A(n175), .Z(n165) );
  GTECH_NAND2 U167 ( .A(I_a[6]), .B(I_b[4]), .Z(n175) );
  GTECH_XOR3 U168 ( .A(n171), .B(n173), .C(n172), .Z(n164) );
  GTECH_OAI21 U169 ( .A(n189), .B(n190), .C(n191), .Z(n172) );
  GTECH_OAI21 U170 ( .A(n192), .B(n193), .C(n194), .Z(n191) );
  GTECH_NOT U171 ( .A(n193), .Z(n189) );
  GTECH_NOT U172 ( .A(n195), .Z(n173) );
  GTECH_NAND2 U173 ( .A(I_b[7]), .B(I_a[3]), .Z(n195) );
  GTECH_NOT U174 ( .A(n169), .Z(n171) );
  GTECH_NAND2 U175 ( .A(I_b[6]), .B(I_a[4]), .Z(n169) );
  GTECH_OAI21 U176 ( .A(n188), .B(n196), .C(n197), .Z(n177) );
  GTECH_OAI21 U177 ( .A(n186), .B(n198), .C(n187), .Z(n197) );
  GTECH_NOT U178 ( .A(n198), .Z(n188) );
  GTECH_NOT U179 ( .A(n199), .Z(n166) );
  GTECH_NAND2 U180 ( .A(I_a[5]), .B(I_b[5]), .Z(n199) );
  GTECH_NOT U181 ( .A(n153), .Z(n157) );
  GTECH_XOR2 U182 ( .A(n179), .B(n150), .Z(n153) );
  GTECH_AOI2N2 U183 ( .A(n200), .B(n201), .C(n202), .D(n203), .Z(n150) );
  GTECH_NAND2 U184 ( .A(n202), .B(n203), .Z(n201) );
  GTECH_XOR2 U185 ( .A(n204), .B(n148), .Z(n179) );
  GTECH_AND2 U186 ( .A(n205), .B(n206), .Z(n148) );
  GTECH_OR_NOT U187 ( .A(n207), .B(n208), .Z(n206) );
  GTECH_OAI21 U188 ( .A(n209), .B(n208), .C(n210), .Z(n205) );
  GTECH_NAND2 U189 ( .A(I_a[7]), .B(I_b[3]), .Z(n204) );
  GTECH_NOT U190 ( .A(n158), .Z(n152) );
  GTECH_OAI2N2 U191 ( .A(n211), .B(n212), .C(n213), .D(n214), .Z(n158) );
  GTECH_NAND2 U192 ( .A(n211), .B(n212), .Z(n214) );
  GTECH_XOR3 U193 ( .A(n211), .B(n215), .C(n216), .Z(N149) );
  GTECH_NOT U194 ( .A(n213), .Z(n216) );
  GTECH_XOR2 U195 ( .A(n217), .B(n182), .Z(n213) );
  GTECH_ADD_ABC U196 ( .A(n218), .B(n219), .C(n220), .COUT(n182) );
  GTECH_XOR3 U197 ( .A(n221), .B(n222), .C(n223), .Z(n219) );
  GTECH_OA21 U198 ( .A(n224), .B(n225), .C(n226), .Z(n218) );
  GTECH_XNOR4 U199 ( .A(n187), .B(n198), .C(n185), .D(n186), .Z(n217) );
  GTECH_NOT U200 ( .A(n196), .Z(n186) );
  GTECH_NAND2 U201 ( .A(I_a[5]), .B(I_b[4]), .Z(n196) );
  GTECH_XOR3 U202 ( .A(n192), .B(n194), .C(n193), .Z(n185) );
  GTECH_OAI21 U203 ( .A(n227), .B(n228), .C(n229), .Z(n193) );
  GTECH_NOT U204 ( .A(n230), .Z(n194) );
  GTECH_NAND2 U205 ( .A(I_b[7]), .B(I_a[2]), .Z(n230) );
  GTECH_NOT U206 ( .A(n190), .Z(n192) );
  GTECH_NAND2 U207 ( .A(I_b[6]), .B(I_a[3]), .Z(n190) );
  GTECH_OAI21 U208 ( .A(n223), .B(n231), .C(n232), .Z(n198) );
  GTECH_OAI21 U209 ( .A(n221), .B(n233), .C(n222), .Z(n232) );
  GTECH_NOT U210 ( .A(n233), .Z(n223) );
  GTECH_NOT U211 ( .A(n234), .Z(n187) );
  GTECH_NAND2 U212 ( .A(I_b[5]), .B(I_a[4]), .Z(n234) );
  GTECH_NOT U213 ( .A(n212), .Z(n215) );
  GTECH_XOR3 U214 ( .A(n235), .B(n202), .C(n200), .Z(n212) );
  GTECH_XOR3 U215 ( .A(n209), .B(n210), .C(n208), .Z(n200) );
  GTECH_OAI21 U216 ( .A(n236), .B(n237), .C(n238), .Z(n208) );
  GTECH_OAI21 U217 ( .A(n239), .B(n240), .C(n241), .Z(n238) );
  GTECH_NOT U218 ( .A(n240), .Z(n236) );
  GTECH_NOT U219 ( .A(n242), .Z(n210) );
  GTECH_NAND2 U220 ( .A(I_a[6]), .B(I_b[3]), .Z(n242) );
  GTECH_NOT U221 ( .A(n207), .Z(n209) );
  GTECH_NAND2 U222 ( .A(I_a[7]), .B(I_b[2]), .Z(n207) );
  GTECH_ADD_ABC U223 ( .A(n243), .B(n244), .C(n245), .COUT(n202) );
  GTECH_XOR2 U224 ( .A(n246), .B(n247), .Z(n244) );
  GTECH_AND2 U225 ( .A(I_a[7]), .B(I_b[1]), .Z(n247) );
  GTECH_NOT U226 ( .A(n203), .Z(n235) );
  GTECH_NAND2 U227 ( .A(I_a[7]), .B(n248), .Z(n203) );
  GTECH_ADD_ABC U228 ( .A(n249), .B(n250), .C(n251), .COUT(n211) );
  GTECH_XOR3 U229 ( .A(n243), .B(n252), .C(n245), .Z(n250) );
  GTECH_NOT U230 ( .A(n253), .Z(n245) );
  GTECH_XOR3 U231 ( .A(n254), .B(n251), .C(n249), .Z(N148) );
  GTECH_ADD_ABC U232 ( .A(n255), .B(n256), .C(n257), .COUT(n249) );
  GTECH_NOT U233 ( .A(n258), .Z(n257) );
  GTECH_XOR3 U234 ( .A(n259), .B(n260), .C(n261), .Z(n256) );
  GTECH_XOR2 U235 ( .A(n262), .B(n263), .Z(n251) );
  GTECH_OA21 U236 ( .A(n224), .B(n225), .C(n226), .Z(n263) );
  GTECH_OAI21 U237 ( .A(n264), .B(n265), .C(n266), .Z(n226) );
  GTECH_NOT U238 ( .A(n224), .Z(n265) );
  GTECH_XNOR4 U239 ( .A(n222), .B(n233), .C(n220), .D(n221), .Z(n262) );
  GTECH_NOT U240 ( .A(n231), .Z(n221) );
  GTECH_NAND2 U241 ( .A(I_b[4]), .B(I_a[4]), .Z(n231) );
  GTECH_XOR3 U242 ( .A(n267), .B(n268), .C(n229), .Z(n220) );
  GTECH_NAND3 U243 ( .A(I_b[6]), .B(I_a[1]), .C(n269), .Z(n229) );
  GTECH_NOT U244 ( .A(n228), .Z(n268) );
  GTECH_NAND2 U245 ( .A(I_b[7]), .B(I_a[1]), .Z(n228) );
  GTECH_NOT U246 ( .A(n227), .Z(n267) );
  GTECH_NAND2 U247 ( .A(I_b[6]), .B(I_a[2]), .Z(n227) );
  GTECH_OAI21 U248 ( .A(n270), .B(n271), .C(n272), .Z(n233) );
  GTECH_OAI21 U249 ( .A(n273), .B(n274), .C(n275), .Z(n272) );
  GTECH_NOT U250 ( .A(n274), .Z(n270) );
  GTECH_NOT U251 ( .A(n276), .Z(n222) );
  GTECH_NAND2 U252 ( .A(I_b[5]), .B(I_a[3]), .Z(n276) );
  GTECH_XOR3 U253 ( .A(n252), .B(n253), .C(n243), .Z(n254) );
  GTECH_ADD_ABC U254 ( .A(n259), .B(n277), .C(n261), .COUT(n243) );
  GTECH_NOT U255 ( .A(n278), .Z(n261) );
  GTECH_XOR3 U256 ( .A(n279), .B(n280), .C(n281), .Z(n277) );
  GTECH_XOR3 U257 ( .A(n239), .B(n241), .C(n240), .Z(n253) );
  GTECH_OAI21 U258 ( .A(n282), .B(n283), .C(n284), .Z(n240) );
  GTECH_OAI21 U259 ( .A(n285), .B(n286), .C(n287), .Z(n284) );
  GTECH_NOT U260 ( .A(n286), .Z(n282) );
  GTECH_NOT U261 ( .A(n288), .Z(n241) );
  GTECH_NAND2 U262 ( .A(I_a[5]), .B(I_b[3]), .Z(n288) );
  GTECH_NOT U263 ( .A(n237), .Z(n239) );
  GTECH_NAND2 U264 ( .A(I_a[6]), .B(I_b[2]), .Z(n237) );
  GTECH_XOR2 U265 ( .A(n289), .B(n246), .Z(n252) );
  GTECH_NOT U266 ( .A(n248), .Z(n246) );
  GTECH_OAI21 U267 ( .A(n281), .B(n290), .C(n291), .Z(n248) );
  GTECH_OAI21 U268 ( .A(n279), .B(n292), .C(n280), .Z(n291) );
  GTECH_NOT U269 ( .A(n292), .Z(n281) );
  GTECH_AND2 U270 ( .A(I_a[7]), .B(I_b[1]), .Z(n289) );
  GTECH_XOR2 U271 ( .A(n293), .B(n255), .Z(N147) );
  GTECH_ADD_ABC U272 ( .A(n294), .B(n295), .C(n296), .COUT(n255) );
  GTECH_XOR3 U273 ( .A(n297), .B(n298), .C(n299), .Z(n295) );
  GTECH_NOT U274 ( .A(n300), .Z(n298) );
  GTECH_OA21 U275 ( .A(n301), .B(n302), .C(n303), .Z(n294) );
  GTECH_XNOR4 U276 ( .A(n260), .B(n278), .C(n258), .D(n259), .Z(n293) );
  GTECH_ADD_ABC U277 ( .A(n297), .B(n304), .C(n299), .COUT(n259) );
  GTECH_NOT U278 ( .A(n305), .Z(n299) );
  GTECH_XOR3 U279 ( .A(n306), .B(n307), .C(n308), .Z(n304) );
  GTECH_XOR3 U280 ( .A(n266), .B(n225), .C(n224), .Z(n258) );
  GTECH_XOR2 U281 ( .A(n309), .B(n269), .Z(n224) );
  GTECH_NOT U282 ( .A(n310), .Z(n269) );
  GTECH_NAND2 U283 ( .A(I_b[7]), .B(I_a[0]), .Z(n310) );
  GTECH_NAND2 U284 ( .A(I_b[6]), .B(I_a[1]), .Z(n309) );
  GTECH_NOT U285 ( .A(n264), .Z(n225) );
  GTECH_XOR3 U286 ( .A(n273), .B(n275), .C(n274), .Z(n264) );
  GTECH_OAI21 U287 ( .A(n311), .B(n312), .C(n313), .Z(n274) );
  GTECH_NOT U288 ( .A(n314), .Z(n275) );
  GTECH_NAND2 U289 ( .A(I_b[5]), .B(I_a[2]), .Z(n314) );
  GTECH_NOT U290 ( .A(n271), .Z(n273) );
  GTECH_NAND2 U291 ( .A(I_b[4]), .B(I_a[3]), .Z(n271) );
  GTECH_NOT U292 ( .A(n315), .Z(n266) );
  GTECH_NAND3 U293 ( .A(I_a[0]), .B(n316), .C(I_b[6]), .Z(n315) );
  GTECH_NOT U294 ( .A(n317), .Z(n316) );
  GTECH_XOR3 U295 ( .A(n285), .B(n287), .C(n286), .Z(n278) );
  GTECH_OAI21 U296 ( .A(n318), .B(n319), .C(n320), .Z(n286) );
  GTECH_OAI21 U297 ( .A(n321), .B(n322), .C(n323), .Z(n320) );
  GTECH_NOT U298 ( .A(n322), .Z(n318) );
  GTECH_NOT U299 ( .A(n324), .Z(n287) );
  GTECH_NAND2 U300 ( .A(I_b[3]), .B(I_a[4]), .Z(n324) );
  GTECH_NOT U301 ( .A(n283), .Z(n285) );
  GTECH_NAND2 U302 ( .A(I_a[5]), .B(I_b[2]), .Z(n283) );
  GTECH_NOT U303 ( .A(n325), .Z(n260) );
  GTECH_XOR3 U304 ( .A(n279), .B(n280), .C(n292), .Z(n325) );
  GTECH_OAI21 U305 ( .A(n308), .B(n326), .C(n327), .Z(n292) );
  GTECH_OAI21 U306 ( .A(n306), .B(n328), .C(n307), .Z(n327) );
  GTECH_NOT U307 ( .A(n328), .Z(n308) );
  GTECH_NOT U308 ( .A(n329), .Z(n280) );
  GTECH_NAND2 U309 ( .A(I_a[6]), .B(I_b[1]), .Z(n329) );
  GTECH_NOT U310 ( .A(n290), .Z(n279) );
  GTECH_NAND2 U311 ( .A(I_a[7]), .B(I_b[0]), .Z(n290) );
  GTECH_XOR2 U312 ( .A(n330), .B(n331), .Z(N146) );
  GTECH_XNOR4 U313 ( .A(n305), .B(n297), .C(n300), .D(n296), .Z(n331) );
  GTECH_XOR2 U314 ( .A(n317), .B(n332), .Z(n296) );
  GTECH_AND2 U315 ( .A(I_b[6]), .B(I_a[0]), .Z(n332) );
  GTECH_XOR3 U316 ( .A(n333), .B(n334), .C(n313), .Z(n317) );
  GTECH_NAND3 U317 ( .A(I_b[4]), .B(I_a[1]), .C(n335), .Z(n313) );
  GTECH_NOT U318 ( .A(n312), .Z(n334) );
  GTECH_NAND2 U319 ( .A(I_b[5]), .B(I_a[1]), .Z(n312) );
  GTECH_NOT U320 ( .A(n311), .Z(n333) );
  GTECH_NAND2 U321 ( .A(I_b[4]), .B(I_a[2]), .Z(n311) );
  GTECH_XOR3 U322 ( .A(n306), .B(n307), .C(n328), .Z(n300) );
  GTECH_OAI21 U323 ( .A(n336), .B(n337), .C(n338), .Z(n328) );
  GTECH_OAI21 U324 ( .A(n339), .B(n340), .C(n341), .Z(n338) );
  GTECH_NOT U325 ( .A(n342), .Z(n307) );
  GTECH_NAND2 U326 ( .A(I_a[5]), .B(I_b[1]), .Z(n342) );
  GTECH_NOT U327 ( .A(n326), .Z(n306) );
  GTECH_NAND2 U328 ( .A(I_a[6]), .B(I_b[0]), .Z(n326) );
  GTECH_ADD_ABC U329 ( .A(n343), .B(n344), .C(n345), .COUT(n297) );
  GTECH_NOT U330 ( .A(n346), .Z(n345) );
  GTECH_XOR3 U331 ( .A(n339), .B(n341), .C(n336), .Z(n344) );
  GTECH_NOT U332 ( .A(n340), .Z(n336) );
  GTECH_XOR3 U333 ( .A(n321), .B(n323), .C(n322), .Z(n305) );
  GTECH_OAI21 U334 ( .A(n347), .B(n348), .C(n349), .Z(n322) );
  GTECH_OAI21 U335 ( .A(n350), .B(n351), .C(n352), .Z(n349) );
  GTECH_NOT U336 ( .A(n351), .Z(n347) );
  GTECH_NOT U337 ( .A(n353), .Z(n323) );
  GTECH_NAND2 U338 ( .A(I_b[3]), .B(I_a[3]), .Z(n353) );
  GTECH_NOT U339 ( .A(n319), .Z(n321) );
  GTECH_NAND2 U340 ( .A(I_b[2]), .B(I_a[4]), .Z(n319) );
  GTECH_OA21 U341 ( .A(n301), .B(n302), .C(n303), .Z(n330) );
  GTECH_OAI21 U342 ( .A(n354), .B(n355), .C(n356), .Z(n303) );
  GTECH_NOT U343 ( .A(n301), .Z(n355) );
  GTECH_XOR3 U344 ( .A(n356), .B(n302), .C(n301), .Z(N145) );
  GTECH_XOR2 U345 ( .A(n357), .B(n335), .Z(n301) );
  GTECH_NOT U346 ( .A(n358), .Z(n335) );
  GTECH_NAND2 U347 ( .A(I_b[5]), .B(I_a[0]), .Z(n358) );
  GTECH_NAND2 U348 ( .A(I_b[4]), .B(I_a[1]), .Z(n357) );
  GTECH_NOT U349 ( .A(n354), .Z(n302) );
  GTECH_XOR2 U350 ( .A(n359), .B(n343), .Z(n354) );
  GTECH_ADD_ABC U351 ( .A(n360), .B(n361), .C(n362), .COUT(n343) );
  GTECH_XOR3 U352 ( .A(n363), .B(n364), .C(n365), .Z(n361) );
  GTECH_OA21 U353 ( .A(n366), .B(n367), .C(n368), .Z(n360) );
  GTECH_XNOR4 U354 ( .A(n341), .B(n340), .C(n346), .D(n339), .Z(n359) );
  GTECH_NOT U355 ( .A(n337), .Z(n339) );
  GTECH_NAND2 U356 ( .A(I_a[5]), .B(I_b[0]), .Z(n337) );
  GTECH_XOR3 U357 ( .A(n350), .B(n352), .C(n351), .Z(n346) );
  GTECH_OAI21 U358 ( .A(n369), .B(n370), .C(n371), .Z(n351) );
  GTECH_NOT U359 ( .A(n372), .Z(n352) );
  GTECH_NAND2 U360 ( .A(I_b[3]), .B(I_a[2]), .Z(n372) );
  GTECH_NOT U361 ( .A(n348), .Z(n350) );
  GTECH_NAND2 U362 ( .A(I_b[2]), .B(I_a[3]), .Z(n348) );
  GTECH_OAI21 U363 ( .A(n365), .B(n373), .C(n374), .Z(n340) );
  GTECH_OAI21 U364 ( .A(n363), .B(n375), .C(n364), .Z(n374) );
  GTECH_NOT U365 ( .A(n373), .Z(n363) );
  GTECH_NOT U366 ( .A(n375), .Z(n365) );
  GTECH_NOT U367 ( .A(n376), .Z(n341) );
  GTECH_NAND2 U368 ( .A(I_a[4]), .B(I_b[1]), .Z(n376) );
  GTECH_NOT U369 ( .A(n377), .Z(n356) );
  GTECH_NAND3 U370 ( .A(I_a[0]), .B(n378), .C(I_b[4]), .Z(n377) );
  GTECH_XOR2 U371 ( .A(n379), .B(n378), .Z(N144) );
  GTECH_XOR2 U372 ( .A(n380), .B(n381), .Z(n378) );
  GTECH_XNOR4 U373 ( .A(n364), .B(n375), .C(n373), .D(n362), .Z(n381) );
  GTECH_XOR3 U374 ( .A(n382), .B(n383), .C(n371), .Z(n362) );
  GTECH_NAND3 U375 ( .A(I_b[2]), .B(I_a[1]), .C(n384), .Z(n371) );
  GTECH_NOT U376 ( .A(n370), .Z(n383) );
  GTECH_NAND2 U377 ( .A(I_b[3]), .B(I_a[1]), .Z(n370) );
  GTECH_NOT U378 ( .A(n369), .Z(n382) );
  GTECH_NAND2 U379 ( .A(I_b[2]), .B(I_a[2]), .Z(n369) );
  GTECH_NAND2 U380 ( .A(I_a[4]), .B(I_b[0]), .Z(n373) );
  GTECH_OAI21 U381 ( .A(n385), .B(n386), .C(n387), .Z(n375) );
  GTECH_OAI21 U382 ( .A(n388), .B(n389), .C(n390), .Z(n387) );
  GTECH_NOT U383 ( .A(n389), .Z(n385) );
  GTECH_NOT U384 ( .A(n391), .Z(n364) );
  GTECH_NAND2 U385 ( .A(I_a[3]), .B(I_b[1]), .Z(n391) );
  GTECH_OA21 U386 ( .A(n366), .B(n367), .C(n368), .Z(n380) );
  GTECH_OAI21 U387 ( .A(n392), .B(n393), .C(n394), .Z(n368) );
  GTECH_NOT U388 ( .A(n366), .Z(n393) );
  GTECH_AND2 U389 ( .A(I_b[4]), .B(I_a[0]), .Z(n379) );
  GTECH_XOR3 U390 ( .A(n394), .B(n367), .C(n366), .Z(N143) );
  GTECH_XOR2 U391 ( .A(n395), .B(n384), .Z(n366) );
  GTECH_NOT U392 ( .A(n396), .Z(n384) );
  GTECH_NAND2 U393 ( .A(I_b[3]), .B(I_a[0]), .Z(n396) );
  GTECH_NAND2 U394 ( .A(I_b[2]), .B(I_a[1]), .Z(n395) );
  GTECH_NOT U395 ( .A(n392), .Z(n367) );
  GTECH_XOR3 U396 ( .A(n388), .B(n390), .C(n389), .Z(n392) );
  GTECH_OAI21 U397 ( .A(n397), .B(n398), .C(n399), .Z(n389) );
  GTECH_NOT U398 ( .A(n400), .Z(n390) );
  GTECH_NAND2 U399 ( .A(I_b[1]), .B(I_a[2]), .Z(n400) );
  GTECH_NOT U400 ( .A(n386), .Z(n388) );
  GTECH_NAND2 U401 ( .A(I_b[0]), .B(I_a[3]), .Z(n386) );
  GTECH_NOT U402 ( .A(n401), .Z(n394) );
  GTECH_NAND3 U403 ( .A(I_a[0]), .B(n402), .C(I_b[2]), .Z(n401) );
  GTECH_XOR2 U404 ( .A(n403), .B(n402), .Z(N142) );
  GTECH_NOT U405 ( .A(n404), .Z(n402) );
  GTECH_XOR3 U406 ( .A(n405), .B(n406), .C(n399), .Z(n404) );
  GTECH_NAND3 U407 ( .A(n407), .B(I_b[0]), .C(I_a[1]), .Z(n399) );
  GTECH_NOT U408 ( .A(n397), .Z(n406) );
  GTECH_NAND2 U409 ( .A(I_a[1]), .B(I_b[1]), .Z(n397) );
  GTECH_NOT U410 ( .A(n398), .Z(n405) );
  GTECH_NAND2 U411 ( .A(I_b[0]), .B(I_a[2]), .Z(n398) );
  GTECH_AND2 U412 ( .A(I_b[2]), .B(I_a[0]), .Z(n403) );
  GTECH_XOR2 U413 ( .A(n407), .B(n408), .Z(N141) );
  GTECH_AND2 U414 ( .A(I_a[1]), .B(I_b[0]), .Z(n408) );
  GTECH_NOT U415 ( .A(n409), .Z(n407) );
  GTECH_NAND2 U416 ( .A(I_a[0]), .B(I_b[1]), .Z(n409) );
  GTECH_AND2 U417 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

