
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI22 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NOT U83 ( .A(n97), .Z(n96) );
  GTECH_AND2 U84 ( .A(n93), .B(n94), .Z(n95) );
  GTECH_XOR2 U85 ( .A(n90), .B(n98), .Z(n86) );
  GTECH_NOT U86 ( .A(n89), .Z(n98) );
  GTECH_OAI22 U87 ( .A(n99), .B(n100), .C(n101), .D(n102), .Z(n89) );
  GTECH_AND2 U88 ( .A(n99), .B(n100), .Z(n101) );
  GTECH_NOT U89 ( .A(n103), .Z(n99) );
  GTECH_NAND2 U90 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U91 ( .A(n104), .Z(n84) );
  GTECH_NAND2 U92 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_XOR2 U93 ( .A(n106), .B(n105), .Z(N153) );
  GTECH_NOT U94 ( .A(n107), .Z(n105) );
  GTECH_XOR3 U95 ( .A(n108), .B(n93), .C(n97), .Z(n107) );
  GTECH_XOR3 U96 ( .A(n109), .B(n110), .C(n103), .Z(n97) );
  GTECH_OAI22 U97 ( .A(n111), .B(n112), .C(n113), .D(n114), .Z(n103) );
  GTECH_AND2 U98 ( .A(n111), .B(n112), .Z(n113) );
  GTECH_NOT U99 ( .A(n115), .Z(n111) );
  GTECH_NOT U100 ( .A(n102), .Z(n110) );
  GTECH_NAND2 U101 ( .A(I_b[7]), .B(I_a[6]), .Z(n102) );
  GTECH_NOT U102 ( .A(n100), .Z(n109) );
  GTECH_NAND2 U103 ( .A(I_a[7]), .B(I_b[6]), .Z(n100) );
  GTECH_ADD_ABC U104 ( .A(n116), .B(n117), .C(n118), .COUT(n93) );
  GTECH_NOT U105 ( .A(n119), .Z(n118) );
  GTECH_XOR2 U106 ( .A(n120), .B(n121), .Z(n117) );
  GTECH_AND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n121) );
  GTECH_NOT U108 ( .A(n94), .Z(n108) );
  GTECH_NAND2 U109 ( .A(I_a[7]), .B(n122), .Z(n94) );
  GTECH_NOT U110 ( .A(n123), .Z(n106) );
  GTECH_NAND2 U111 ( .A(n124), .B(n125), .Z(n123) );
  GTECH_NOT U112 ( .A(n126), .Z(n125) );
  GTECH_XOR2 U113 ( .A(n126), .B(n127), .Z(N152) );
  GTECH_NOT U114 ( .A(n124), .Z(n127) );
  GTECH_XOR4 U115 ( .A(n128), .B(n120), .C(n116), .D(n119), .Z(n124) );
  GTECH_XOR3 U116 ( .A(n129), .B(n130), .C(n115), .Z(n119) );
  GTECH_OAI22 U117 ( .A(n131), .B(n132), .C(n133), .D(n134), .Z(n115) );
  GTECH_AND2 U118 ( .A(n131), .B(n132), .Z(n133) );
  GTECH_NOT U119 ( .A(n135), .Z(n131) );
  GTECH_NOT U120 ( .A(n114), .Z(n130) );
  GTECH_NAND2 U121 ( .A(I_b[7]), .B(I_a[5]), .Z(n114) );
  GTECH_NOT U122 ( .A(n112), .Z(n129) );
  GTECH_NAND2 U123 ( .A(I_b[6]), .B(I_a[6]), .Z(n112) );
  GTECH_ADD_ABC U124 ( .A(n136), .B(n137), .C(n138), .COUT(n116) );
  GTECH_NOT U125 ( .A(n139), .Z(n138) );
  GTECH_XOR3 U126 ( .A(n140), .B(n141), .C(n142), .Z(n137) );
  GTECH_NOT U127 ( .A(n143), .Z(n140) );
  GTECH_NOT U128 ( .A(n122), .Z(n120) );
  GTECH_OAI22 U129 ( .A(n142), .B(n143), .C(n144), .D(n145), .Z(n122) );
  GTECH_AND2 U130 ( .A(n142), .B(n143), .Z(n144) );
  GTECH_NOT U131 ( .A(n146), .Z(n142) );
  GTECH_AND2 U132 ( .A(I_a[7]), .B(I_b[5]), .Z(n128) );
  GTECH_ADD_ABC U133 ( .A(n147), .B(n148), .C(n149), .COUT(n126) );
  GTECH_NOT U134 ( .A(n150), .Z(n149) );
  GTECH_OA22 U135 ( .A(n151), .B(n152), .C(n153), .D(n154), .Z(n148) );
  GTECH_OA21 U136 ( .A(n155), .B(n156), .C(n157), .Z(n147) );
  GTECH_AO21 U137 ( .A(n155), .B(n156), .C(n158), .Z(n157) );
  GTECH_XOR3 U138 ( .A(n159), .B(n150), .C(n160), .Z(N151) );
  GTECH_OA21 U139 ( .A(n155), .B(n156), .C(n161), .Z(n160) );
  GTECH_AO21 U140 ( .A(n155), .B(n156), .C(n158), .Z(n161) );
  GTECH_XOR2 U141 ( .A(n162), .B(n136), .Z(n150) );
  GTECH_ADD_ABC U142 ( .A(n163), .B(n164), .C(n165), .COUT(n136) );
  GTECH_NOT U143 ( .A(n166), .Z(n165) );
  GTECH_XOR3 U144 ( .A(n167), .B(n168), .C(n169), .Z(n164) );
  GTECH_XOR4 U145 ( .A(n141), .B(n146), .C(n143), .D(n139), .Z(n162) );
  GTECH_XOR3 U146 ( .A(n170), .B(n171), .C(n135), .Z(n139) );
  GTECH_OAI22 U147 ( .A(n172), .B(n173), .C(n174), .D(n175), .Z(n135) );
  GTECH_AND2 U148 ( .A(n172), .B(n173), .Z(n174) );
  GTECH_NOT U149 ( .A(n176), .Z(n172) );
  GTECH_NOT U150 ( .A(n134), .Z(n171) );
  GTECH_NAND2 U151 ( .A(I_b[7]), .B(I_a[4]), .Z(n134) );
  GTECH_NOT U152 ( .A(n132), .Z(n170) );
  GTECH_NAND2 U153 ( .A(I_b[6]), .B(I_a[5]), .Z(n132) );
  GTECH_NAND2 U154 ( .A(I_a[7]), .B(I_b[4]), .Z(n143) );
  GTECH_OAI22 U155 ( .A(n169), .B(n177), .C(n178), .D(n179), .Z(n146) );
  GTECH_AND2 U156 ( .A(n169), .B(n177), .Z(n178) );
  GTECH_NOT U157 ( .A(n180), .Z(n169) );
  GTECH_NOT U158 ( .A(n145), .Z(n141) );
  GTECH_NAND2 U159 ( .A(I_a[6]), .B(I_b[5]), .Z(n145) );
  GTECH_OA22 U160 ( .A(n151), .B(n152), .C(n153), .D(n154), .Z(n159) );
  GTECH_NOT U161 ( .A(n181), .Z(n154) );
  GTECH_NOT U162 ( .A(I_a[7]), .Z(n152) );
  GTECH_XOR3 U163 ( .A(n155), .B(n182), .C(n158), .Z(N150) );
  GTECH_XOR2 U164 ( .A(n163), .B(n183), .Z(n158) );
  GTECH_XOR4 U165 ( .A(n168), .B(n180), .C(n166), .D(n167), .Z(n183) );
  GTECH_NOT U166 ( .A(n177), .Z(n167) );
  GTECH_NAND2 U167 ( .A(I_a[6]), .B(I_b[4]), .Z(n177) );
  GTECH_XOR3 U168 ( .A(n184), .B(n185), .C(n176), .Z(n166) );
  GTECH_OAI22 U169 ( .A(n186), .B(n187), .C(n188), .D(n189), .Z(n176) );
  GTECH_AND2 U170 ( .A(n186), .B(n187), .Z(n188) );
  GTECH_NOT U171 ( .A(n190), .Z(n186) );
  GTECH_NOT U172 ( .A(n175), .Z(n185) );
  GTECH_NAND2 U173 ( .A(I_b[7]), .B(I_a[3]), .Z(n175) );
  GTECH_NOT U174 ( .A(n173), .Z(n184) );
  GTECH_NAND2 U175 ( .A(I_b[6]), .B(I_a[4]), .Z(n173) );
  GTECH_OAI22 U176 ( .A(n191), .B(n192), .C(n193), .D(n194), .Z(n180) );
  GTECH_AND2 U177 ( .A(n191), .B(n192), .Z(n193) );
  GTECH_NOT U178 ( .A(n179), .Z(n168) );
  GTECH_NAND2 U179 ( .A(I_a[5]), .B(I_b[5]), .Z(n179) );
  GTECH_ADD_ABC U180 ( .A(n195), .B(n196), .C(n197), .COUT(n163) );
  GTECH_NOT U181 ( .A(n198), .Z(n197) );
  GTECH_XOR3 U182 ( .A(n199), .B(n200), .C(n191), .Z(n196) );
  GTECH_NOT U183 ( .A(n201), .Z(n191) );
  GTECH_NOT U184 ( .A(n156), .Z(n182) );
  GTECH_XOR2 U185 ( .A(n181), .B(n153), .Z(n156) );
  GTECH_AOI2N2 U186 ( .A(n202), .B(n203), .C(n204), .D(n205), .Z(n153) );
  GTECH_NAND2 U187 ( .A(n204), .B(n205), .Z(n203) );
  GTECH_XOR2 U188 ( .A(n206), .B(n151), .Z(n181) );
  GTECH_OA21 U189 ( .A(n207), .B(n208), .C(n209), .Z(n151) );
  GTECH_AO21 U190 ( .A(n207), .B(n208), .C(n210), .Z(n209) );
  GTECH_NOT U191 ( .A(n211), .Z(n207) );
  GTECH_NAND2 U192 ( .A(I_a[7]), .B(I_b[3]), .Z(n206) );
  GTECH_OA21 U193 ( .A(n212), .B(n213), .C(n214), .Z(n155) );
  GTECH_AO21 U194 ( .A(n212), .B(n213), .C(n215), .Z(n214) );
  GTECH_XOR3 U195 ( .A(n212), .B(n216), .C(n215), .Z(N149) );
  GTECH_XOR2 U196 ( .A(n195), .B(n217), .Z(n215) );
  GTECH_XOR4 U197 ( .A(n200), .B(n201), .C(n198), .D(n199), .Z(n217) );
  GTECH_NOT U198 ( .A(n192), .Z(n199) );
  GTECH_NAND2 U199 ( .A(I_a[5]), .B(I_b[4]), .Z(n192) );
  GTECH_XOR3 U200 ( .A(n218), .B(n219), .C(n190), .Z(n198) );
  GTECH_AO21 U201 ( .A(n220), .B(n221), .C(n222), .Z(n190) );
  GTECH_NOT U202 ( .A(n223), .Z(n222) );
  GTECH_NOT U203 ( .A(n189), .Z(n219) );
  GTECH_NAND2 U204 ( .A(I_b[7]), .B(I_a[2]), .Z(n189) );
  GTECH_NOT U205 ( .A(n187), .Z(n218) );
  GTECH_NAND2 U206 ( .A(I_b[6]), .B(I_a[3]), .Z(n187) );
  GTECH_OAI22 U207 ( .A(n224), .B(n225), .C(n226), .D(n227), .Z(n201) );
  GTECH_AND2 U208 ( .A(n224), .B(n225), .Z(n226) );
  GTECH_NOT U209 ( .A(n194), .Z(n200) );
  GTECH_NAND2 U210 ( .A(I_b[5]), .B(I_a[4]), .Z(n194) );
  GTECH_ADD_ABC U211 ( .A(n228), .B(n229), .C(n230), .COUT(n195) );
  GTECH_XOR3 U212 ( .A(n231), .B(n232), .C(n224), .Z(n229) );
  GTECH_NOT U213 ( .A(n233), .Z(n224) );
  GTECH_NOT U214 ( .A(n225), .Z(n231) );
  GTECH_OA21 U215 ( .A(n234), .B(n235), .C(n236), .Z(n228) );
  GTECH_AO21 U216 ( .A(n234), .B(n235), .C(n237), .Z(n236) );
  GTECH_NOT U217 ( .A(n213), .Z(n216) );
  GTECH_XOR3 U218 ( .A(n238), .B(n204), .C(n202), .Z(n213) );
  GTECH_XOR3 U219 ( .A(n239), .B(n240), .C(n211), .Z(n202) );
  GTECH_OAI22 U220 ( .A(n241), .B(n242), .C(n243), .D(n244), .Z(n211) );
  GTECH_AND2 U221 ( .A(n241), .B(n242), .Z(n243) );
  GTECH_NOT U222 ( .A(n245), .Z(n241) );
  GTECH_NOT U223 ( .A(n210), .Z(n240) );
  GTECH_NAND2 U224 ( .A(I_a[6]), .B(I_b[3]), .Z(n210) );
  GTECH_NOT U225 ( .A(n208), .Z(n239) );
  GTECH_NAND2 U226 ( .A(I_a[7]), .B(I_b[2]), .Z(n208) );
  GTECH_ADD_ABC U227 ( .A(n246), .B(n247), .C(n248), .COUT(n204) );
  GTECH_XOR2 U228 ( .A(n249), .B(n250), .Z(n247) );
  GTECH_AND2 U229 ( .A(I_a[7]), .B(I_b[1]), .Z(n250) );
  GTECH_NOT U230 ( .A(n205), .Z(n238) );
  GTECH_NAND2 U231 ( .A(I_a[7]), .B(n251), .Z(n205) );
  GTECH_ADD_ABC U232 ( .A(n252), .B(n253), .C(n254), .COUT(n212) );
  GTECH_XOR3 U233 ( .A(n246), .B(n255), .C(n248), .Z(n253) );
  GTECH_NOT U234 ( .A(n256), .Z(n248) );
  GTECH_XOR2 U235 ( .A(n252), .B(n257), .Z(N148) );
  GTECH_XOR4 U236 ( .A(n255), .B(n256), .C(n254), .D(n246), .Z(n257) );
  GTECH_ADD_ABC U237 ( .A(n258), .B(n259), .C(n260), .COUT(n246) );
  GTECH_XOR3 U238 ( .A(n261), .B(n262), .C(n263), .Z(n259) );
  GTECH_XOR2 U239 ( .A(n264), .B(n265), .Z(n254) );
  GTECH_OA21 U240 ( .A(n234), .B(n235), .C(n266), .Z(n265) );
  GTECH_AO21 U241 ( .A(n234), .B(n235), .C(n237), .Z(n266) );
  GTECH_XOR4 U242 ( .A(n232), .B(n233), .C(n225), .D(n230), .Z(n264) );
  GTECH_XOR3 U243 ( .A(n221), .B(n220), .C(n223), .Z(n230) );
  GTECH_NAND3 U244 ( .A(I_b[6]), .B(I_a[1]), .C(n267), .Z(n223) );
  GTECH_NOT U245 ( .A(n268), .Z(n220) );
  GTECH_NAND2 U246 ( .A(I_b[7]), .B(I_a[1]), .Z(n268) );
  GTECH_NOT U247 ( .A(n269), .Z(n221) );
  GTECH_NAND2 U248 ( .A(I_b[6]), .B(I_a[2]), .Z(n269) );
  GTECH_NAND2 U249 ( .A(I_b[4]), .B(I_a[4]), .Z(n225) );
  GTECH_OAI22 U250 ( .A(n270), .B(n271), .C(n272), .D(n273), .Z(n233) );
  GTECH_AND2 U251 ( .A(n270), .B(n271), .Z(n272) );
  GTECH_NOT U252 ( .A(n274), .Z(n270) );
  GTECH_NOT U253 ( .A(n227), .Z(n232) );
  GTECH_NAND2 U254 ( .A(I_b[5]), .B(I_a[3]), .Z(n227) );
  GTECH_XOR3 U255 ( .A(n275), .B(n276), .C(n245), .Z(n256) );
  GTECH_OAI22 U256 ( .A(n277), .B(n278), .C(n279), .D(n280), .Z(n245) );
  GTECH_AND2 U257 ( .A(n277), .B(n278), .Z(n279) );
  GTECH_NOT U258 ( .A(n281), .Z(n277) );
  GTECH_NOT U259 ( .A(n244), .Z(n276) );
  GTECH_NAND2 U260 ( .A(I_a[5]), .B(I_b[3]), .Z(n244) );
  GTECH_NOT U261 ( .A(n242), .Z(n275) );
  GTECH_NAND2 U262 ( .A(I_a[6]), .B(I_b[2]), .Z(n242) );
  GTECH_XOR2 U263 ( .A(n282), .B(n249), .Z(n255) );
  GTECH_NOT U264 ( .A(n251), .Z(n249) );
  GTECH_OAI22 U265 ( .A(n263), .B(n283), .C(n284), .D(n285), .Z(n251) );
  GTECH_AND2 U266 ( .A(n263), .B(n283), .Z(n284) );
  GTECH_NOT U267 ( .A(n286), .Z(n263) );
  GTECH_AND2 U268 ( .A(I_a[7]), .B(I_b[1]), .Z(n282) );
  GTECH_ADD_ABC U269 ( .A(n287), .B(n288), .C(n289), .COUT(n252) );
  GTECH_NOT U270 ( .A(n290), .Z(n289) );
  GTECH_XOR3 U271 ( .A(n258), .B(n291), .C(n260), .Z(n288) );
  GTECH_NOT U272 ( .A(n292), .Z(n260) );
  GTECH_NOT U273 ( .A(n293), .Z(n291) );
  GTECH_XOR2 U274 ( .A(n294), .B(n287), .Z(N147) );
  GTECH_ADD_ABC U275 ( .A(n295), .B(n296), .C(n297), .COUT(n287) );
  GTECH_XOR3 U276 ( .A(n298), .B(n299), .C(n300), .Z(n296) );
  GTECH_OA21 U277 ( .A(n301), .B(n302), .C(n303), .Z(n295) );
  GTECH_AO21 U278 ( .A(n301), .B(n302), .C(n304), .Z(n303) );
  GTECH_XOR4 U279 ( .A(n292), .B(n258), .C(n293), .D(n290), .Z(n294) );
  GTECH_XOR3 U280 ( .A(n305), .B(n235), .C(n234), .Z(n290) );
  GTECH_XOR2 U281 ( .A(n306), .B(n267), .Z(n234) );
  GTECH_NOT U282 ( .A(n307), .Z(n267) );
  GTECH_NAND2 U283 ( .A(I_b[7]), .B(I_a[0]), .Z(n307) );
  GTECH_NAND2 U284 ( .A(I_b[6]), .B(I_a[1]), .Z(n306) );
  GTECH_NOT U285 ( .A(n308), .Z(n235) );
  GTECH_XOR3 U286 ( .A(n309), .B(n310), .C(n274), .Z(n308) );
  GTECH_AO21 U287 ( .A(n311), .B(n312), .C(n313), .Z(n274) );
  GTECH_NOT U288 ( .A(n314), .Z(n313) );
  GTECH_NOT U289 ( .A(n273), .Z(n310) );
  GTECH_NAND2 U290 ( .A(I_b[5]), .B(I_a[2]), .Z(n273) );
  GTECH_NOT U291 ( .A(n271), .Z(n309) );
  GTECH_NAND2 U292 ( .A(I_b[4]), .B(I_a[3]), .Z(n271) );
  GTECH_NOT U293 ( .A(n237), .Z(n305) );
  GTECH_NAND3 U294 ( .A(I_a[0]), .B(n315), .C(I_b[6]), .Z(n237) );
  GTECH_NOT U295 ( .A(n316), .Z(n315) );
  GTECH_XOR3 U296 ( .A(n261), .B(n262), .C(n286), .Z(n293) );
  GTECH_OAI22 U297 ( .A(n317), .B(n318), .C(n319), .D(n320), .Z(n286) );
  GTECH_AND2 U298 ( .A(n317), .B(n318), .Z(n319) );
  GTECH_NOT U299 ( .A(n285), .Z(n262) );
  GTECH_NAND2 U300 ( .A(I_a[6]), .B(I_b[1]), .Z(n285) );
  GTECH_NOT U301 ( .A(n283), .Z(n261) );
  GTECH_NAND2 U302 ( .A(I_a[7]), .B(I_b[0]), .Z(n283) );
  GTECH_ADD_ABC U303 ( .A(n298), .B(n321), .C(n300), .COUT(n258) );
  GTECH_NOT U304 ( .A(n322), .Z(n300) );
  GTECH_XOR3 U305 ( .A(n323), .B(n324), .C(n317), .Z(n321) );
  GTECH_NOT U306 ( .A(n325), .Z(n317) );
  GTECH_XOR3 U307 ( .A(n326), .B(n327), .C(n281), .Z(n292) );
  GTECH_OAI22 U308 ( .A(n328), .B(n329), .C(n330), .D(n331), .Z(n281) );
  GTECH_AND2 U309 ( .A(n328), .B(n329), .Z(n330) );
  GTECH_NOT U310 ( .A(n332), .Z(n328) );
  GTECH_NOT U311 ( .A(n280), .Z(n327) );
  GTECH_NAND2 U312 ( .A(I_b[3]), .B(I_a[4]), .Z(n280) );
  GTECH_NOT U313 ( .A(n278), .Z(n326) );
  GTECH_NAND2 U314 ( .A(I_a[5]), .B(I_b[2]), .Z(n278) );
  GTECH_XOR2 U315 ( .A(n333), .B(n334), .Z(N146) );
  GTECH_XOR4 U316 ( .A(n299), .B(n322), .C(n297), .D(n298), .Z(n334) );
  GTECH_ADD_ABC U317 ( .A(n335), .B(n336), .C(n337), .COUT(n298) );
  GTECH_NOT U318 ( .A(n338), .Z(n337) );
  GTECH_XOR3 U319 ( .A(n339), .B(n340), .C(n341), .Z(n336) );
  GTECH_XOR2 U320 ( .A(n316), .B(n342), .Z(n297) );
  GTECH_AND2 U321 ( .A(I_b[6]), .B(I_a[0]), .Z(n342) );
  GTECH_XOR3 U322 ( .A(n312), .B(n311), .C(n314), .Z(n316) );
  GTECH_NAND3 U323 ( .A(I_b[4]), .B(I_a[1]), .C(n343), .Z(n314) );
  GTECH_NOT U324 ( .A(n344), .Z(n311) );
  GTECH_NAND2 U325 ( .A(I_b[5]), .B(I_a[1]), .Z(n344) );
  GTECH_NOT U326 ( .A(n345), .Z(n312) );
  GTECH_NAND2 U327 ( .A(I_b[4]), .B(I_a[2]), .Z(n345) );
  GTECH_XOR3 U328 ( .A(n346), .B(n347), .C(n332), .Z(n322) );
  GTECH_OAI22 U329 ( .A(n348), .B(n349), .C(n350), .D(n351), .Z(n332) );
  GTECH_AND2 U330 ( .A(n348), .B(n349), .Z(n350) );
  GTECH_NOT U331 ( .A(n352), .Z(n348) );
  GTECH_NOT U332 ( .A(n331), .Z(n347) );
  GTECH_NAND2 U333 ( .A(I_b[3]), .B(I_a[3]), .Z(n331) );
  GTECH_NOT U334 ( .A(n329), .Z(n346) );
  GTECH_NAND2 U335 ( .A(I_b[2]), .B(I_a[4]), .Z(n329) );
  GTECH_NOT U336 ( .A(n353), .Z(n299) );
  GTECH_XOR3 U337 ( .A(n323), .B(n324), .C(n325), .Z(n353) );
  GTECH_OAI22 U338 ( .A(n341), .B(n354), .C(n355), .D(n356), .Z(n325) );
  GTECH_AND2 U339 ( .A(n341), .B(n354), .Z(n355) );
  GTECH_NOT U340 ( .A(n357), .Z(n341) );
  GTECH_NOT U341 ( .A(n320), .Z(n324) );
  GTECH_NAND2 U342 ( .A(I_a[5]), .B(I_b[1]), .Z(n320) );
  GTECH_NOT U343 ( .A(n318), .Z(n323) );
  GTECH_NAND2 U344 ( .A(I_a[6]), .B(I_b[0]), .Z(n318) );
  GTECH_OA21 U345 ( .A(n301), .B(n302), .C(n358), .Z(n333) );
  GTECH_AO21 U346 ( .A(n301), .B(n302), .C(n304), .Z(n358) );
  GTECH_XOR3 U347 ( .A(n359), .B(n302), .C(n301), .Z(N145) );
  GTECH_XOR2 U348 ( .A(n360), .B(n343), .Z(n301) );
  GTECH_NOT U349 ( .A(n361), .Z(n343) );
  GTECH_NAND2 U350 ( .A(I_b[5]), .B(I_a[0]), .Z(n361) );
  GTECH_NAND2 U351 ( .A(I_b[4]), .B(I_a[1]), .Z(n360) );
  GTECH_XOR2 U352 ( .A(n335), .B(n362), .Z(n302) );
  GTECH_XOR4 U353 ( .A(n340), .B(n357), .C(n338), .D(n339), .Z(n362) );
  GTECH_NOT U354 ( .A(n354), .Z(n339) );
  GTECH_NAND2 U355 ( .A(I_a[5]), .B(I_b[0]), .Z(n354) );
  GTECH_XOR3 U356 ( .A(n363), .B(n364), .C(n352), .Z(n338) );
  GTECH_AO21 U357 ( .A(n365), .B(n366), .C(n367), .Z(n352) );
  GTECH_NOT U358 ( .A(n368), .Z(n367) );
  GTECH_NOT U359 ( .A(n351), .Z(n364) );
  GTECH_NAND2 U360 ( .A(I_b[3]), .B(I_a[2]), .Z(n351) );
  GTECH_NOT U361 ( .A(n349), .Z(n363) );
  GTECH_NAND2 U362 ( .A(I_b[2]), .B(I_a[3]), .Z(n349) );
  GTECH_OAI22 U363 ( .A(n369), .B(n370), .C(n371), .D(n372), .Z(n357) );
  GTECH_AND2 U364 ( .A(n369), .B(n370), .Z(n371) );
  GTECH_NOT U365 ( .A(n356), .Z(n340) );
  GTECH_NAND2 U366 ( .A(I_a[4]), .B(I_b[1]), .Z(n356) );
  GTECH_ADD_ABC U367 ( .A(n373), .B(n374), .C(n375), .COUT(n335) );
  GTECH_XOR3 U368 ( .A(n376), .B(n377), .C(n369), .Z(n374) );
  GTECH_NOT U369 ( .A(n378), .Z(n369) );
  GTECH_OA21 U370 ( .A(n379), .B(n380), .C(n381), .Z(n373) );
  GTECH_AO21 U371 ( .A(n379), .B(n380), .C(n382), .Z(n381) );
  GTECH_NOT U372 ( .A(n304), .Z(n359) );
  GTECH_NAND3 U373 ( .A(I_a[0]), .B(n383), .C(I_b[4]), .Z(n304) );
  GTECH_XOR2 U374 ( .A(n384), .B(n383), .Z(N144) );
  GTECH_XOR2 U375 ( .A(n385), .B(n386), .Z(n383) );
  GTECH_XOR4 U376 ( .A(n377), .B(n378), .C(n375), .D(n376), .Z(n386) );
  GTECH_NOT U377 ( .A(n370), .Z(n376) );
  GTECH_NAND2 U378 ( .A(I_a[4]), .B(I_b[0]), .Z(n370) );
  GTECH_XOR3 U379 ( .A(n366), .B(n365), .C(n368), .Z(n375) );
  GTECH_NAND3 U380 ( .A(I_b[2]), .B(I_a[1]), .C(n387), .Z(n368) );
  GTECH_NOT U381 ( .A(n388), .Z(n365) );
  GTECH_NAND2 U382 ( .A(I_b[3]), .B(I_a[1]), .Z(n388) );
  GTECH_NOT U383 ( .A(n389), .Z(n366) );
  GTECH_NAND2 U384 ( .A(I_b[2]), .B(I_a[2]), .Z(n389) );
  GTECH_OAI22 U385 ( .A(n390), .B(n391), .C(n392), .D(n393), .Z(n378) );
  GTECH_AND2 U386 ( .A(n390), .B(n391), .Z(n392) );
  GTECH_NOT U387 ( .A(n394), .Z(n390) );
  GTECH_NOT U388 ( .A(n372), .Z(n377) );
  GTECH_NAND2 U389 ( .A(I_a[3]), .B(I_b[1]), .Z(n372) );
  GTECH_OA21 U390 ( .A(n379), .B(n380), .C(n395), .Z(n385) );
  GTECH_AO21 U391 ( .A(n379), .B(n380), .C(n382), .Z(n395) );
  GTECH_AND2 U392 ( .A(I_b[4]), .B(I_a[0]), .Z(n384) );
  GTECH_XOR3 U393 ( .A(n396), .B(n380), .C(n379), .Z(N143) );
  GTECH_XOR2 U394 ( .A(n397), .B(n387), .Z(n379) );
  GTECH_NOT U395 ( .A(n398), .Z(n387) );
  GTECH_NAND2 U396 ( .A(I_b[3]), .B(I_a[0]), .Z(n398) );
  GTECH_NAND2 U397 ( .A(I_b[2]), .B(I_a[1]), .Z(n397) );
  GTECH_NOT U398 ( .A(n399), .Z(n380) );
  GTECH_XOR3 U399 ( .A(n400), .B(n401), .C(n394), .Z(n399) );
  GTECH_AO21 U400 ( .A(n402), .B(n403), .C(n404), .Z(n394) );
  GTECH_NOT U401 ( .A(n405), .Z(n404) );
  GTECH_NOT U402 ( .A(n393), .Z(n401) );
  GTECH_NAND2 U403 ( .A(I_b[1]), .B(I_a[2]), .Z(n393) );
  GTECH_NOT U404 ( .A(n391), .Z(n400) );
  GTECH_NAND2 U405 ( .A(I_b[0]), .B(I_a[3]), .Z(n391) );
  GTECH_NOT U406 ( .A(n382), .Z(n396) );
  GTECH_NAND3 U407 ( .A(I_a[0]), .B(n406), .C(I_b[2]), .Z(n382) );
  GTECH_XOR2 U408 ( .A(n407), .B(n406), .Z(N142) );
  GTECH_NOT U409 ( .A(n408), .Z(n406) );
  GTECH_XOR3 U410 ( .A(n402), .B(n403), .C(n405), .Z(n408) );
  GTECH_NAND3 U411 ( .A(n409), .B(I_b[0]), .C(I_a[1]), .Z(n405) );
  GTECH_NOT U412 ( .A(n410), .Z(n403) );
  GTECH_NAND2 U413 ( .A(I_a[1]), .B(I_b[1]), .Z(n410) );
  GTECH_NOT U414 ( .A(n411), .Z(n402) );
  GTECH_NAND2 U415 ( .A(I_b[0]), .B(I_a[2]), .Z(n411) );
  GTECH_AND2 U416 ( .A(I_b[2]), .B(I_a[0]), .Z(n407) );
  GTECH_XOR2 U417 ( .A(n409), .B(n412), .Z(N141) );
  GTECH_AND2 U418 ( .A(I_a[1]), .B(I_b[0]), .Z(n412) );
  GTECH_NOT U419 ( .A(n413), .Z(n409) );
  GTECH_NAND2 U420 ( .A(I_a[0]), .B(I_b[1]), .Z(n413) );
  GTECH_AND2 U421 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

