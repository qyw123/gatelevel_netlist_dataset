
module bcd_counter ( clk, reset, ena, q );
  output [3:1] ena;
  output [15:0] q;
  input clk, reset;
  wire   N10, N11, N12, N13, N22, N23, N24, N25, N26, N38, N39, N40, N41, N42,
         N54, N55, N56, N57, N58, n50, n62, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130;

  GTECH_FD2 ones_reg_0_ ( .D(N10), .CP(clk), .CD(n62), .Q(q[0]) );
  GTECH_FD2 ones_reg_2_ ( .D(N12), .CP(clk), .CD(n62), .Q(q[2]) );
  GTECH_FD2 ones_reg_1_ ( .D(N11), .CP(clk), .CD(n62), .Q(q[1]) );
  GTECH_FD2 ones_reg_3_ ( .D(N13), .CP(clk), .CD(n62), .Q(q[3]) );
  GTECH_FJK1S tens_reg_0_ ( .J(n50), .K(n50), .TI(N22), .TE(N25), .CP(clk), 
        .Q(q[4]) );
  GTECH_FJK1S tens_reg_2_ ( .J(n50), .K(n50), .TI(N24), .TE(N25), .CP(clk), 
        .Q(q[6]) );
  GTECH_FJK1S tens_reg_1_ ( .J(n50), .K(n50), .TI(N23), .TE(N25), .CP(clk), 
        .Q(q[5]) );
  GTECH_FJK1S tens_reg_3_ ( .J(n50), .K(n50), .TI(N26), .TE(N25), .CP(clk), 
        .Q(q[7]) );
  GTECH_FJK1S hundreds_reg_0_ ( .J(n50), .K(n50), .TI(N38), .TE(N41), .CP(clk), 
        .Q(q[8]) );
  GTECH_FJK1S hundreds_reg_2_ ( .J(n50), .K(n50), .TI(N40), .TE(N41), .CP(clk), 
        .Q(q[10]) );
  GTECH_FJK1S hundreds_reg_1_ ( .J(n50), .K(n50), .TI(N39), .TE(N41), .CP(clk), 
        .Q(q[9]) );
  GTECH_FJK1S hundreds_reg_3_ ( .J(n50), .K(n50), .TI(N42), .TE(N41), .CP(clk), 
        .Q(q[11]) );
  GTECH_FJK1S thousands_reg_0_ ( .J(n50), .K(n50), .TI(N54), .TE(N57), .CP(clk), .Q(q[12]) );
  GTECH_FJK1S thousands_reg_2_ ( .J(n50), .K(n50), .TI(N56), .TE(N57), .CP(clk), .Q(q[14]) );
  GTECH_FJK1S thousands_reg_1_ ( .J(n50), .K(n50), .TI(N55), .TE(N57), .CP(clk), .Q(q[13]) );
  GTECH_FJK1S thousands_reg_3_ ( .J(n50), .K(n50), .TI(N58), .TE(N57), .CP(clk), .Q(q[15]) );
  GTECH_ONE U85 ( .Z(n62) );
  GTECH_ZERO U86 ( .Z(n50) );
  GTECH_MUX2 U87 ( .A(n78), .B(n79), .S(q[15]), .Z(N58) );
  GTECH_AO21 U88 ( .A(n80), .B(n81), .C(n82), .Z(n79) );
  GTECH_AND2 U89 ( .A(q[14]), .B(n83), .Z(n78) );
  GTECH_MUX2 U90 ( .A(n83), .B(n82), .S(q[14]), .Z(N56) );
  GTECH_AO21 U91 ( .A(n80), .B(n84), .C(N54), .Z(n82) );
  GTECH_NOT U92 ( .A(n85), .Z(n83) );
  GTECH_NAND3 U93 ( .A(n80), .B(q[12]), .C(q[13]), .Z(n85) );
  GTECH_MUX2 U94 ( .A(n86), .B(N54), .S(q[13]), .Z(N55) );
  GTECH_AND2 U95 ( .A(n80), .B(q[12]), .Z(n86) );
  GTECH_NOT U96 ( .A(n87), .Z(N54) );
  GTECH_NAND2 U97 ( .A(n80), .B(n88), .Z(n87) );
  GTECH_NOT U98 ( .A(q[12]), .Z(n88) );
  GTECH_AND3 U99 ( .A(n89), .B(ena[3]), .C(n90), .Z(n80) );
  GTECH_NAND4 U100 ( .A(q[15]), .B(q[12]), .C(n84), .D(n81), .Z(n90) );
  GTECH_NOT U101 ( .A(q[14]), .Z(n81) );
  GTECH_NOT U102 ( .A(q[13]), .Z(n84) );
  GTECH_NOT U103 ( .A(n91), .Z(ena[3]) );
  GTECH_MUX2 U104 ( .A(n92), .B(n93), .S(q[11]), .Z(N42) );
  GTECH_AO21 U105 ( .A(n94), .B(n95), .C(n96), .Z(n93) );
  GTECH_AND2 U106 ( .A(q[10]), .B(n97), .Z(n92) );
  GTECH_NAND2 U107 ( .A(n98), .B(n99), .Z(N41) );
  GTECH_MUX2 U108 ( .A(n97), .B(n96), .S(q[10]), .Z(N40) );
  GTECH_AO21 U109 ( .A(n94), .B(n100), .C(N38), .Z(n96) );
  GTECH_NOT U110 ( .A(n101), .Z(n97) );
  GTECH_NAND3 U111 ( .A(n94), .B(q[8]), .C(q[9]), .Z(n101) );
  GTECH_MUX2 U112 ( .A(n102), .B(N38), .S(q[9]), .Z(N39) );
  GTECH_AND2 U113 ( .A(n94), .B(q[8]), .Z(n102) );
  GTECH_NOT U114 ( .A(n103), .Z(N38) );
  GTECH_NAND2 U115 ( .A(n94), .B(n104), .Z(n103) );
  GTECH_NOT U116 ( .A(q[8]), .Z(n104) );
  GTECH_NOT U117 ( .A(n98), .Z(n94) );
  GTECH_NAND2 U118 ( .A(ena[2]), .B(n99), .Z(n98) );
  GTECH_NOT U119 ( .A(N57), .Z(n99) );
  GTECH_NAND2 U120 ( .A(n89), .B(n91), .Z(N57) );
  GTECH_NAND5 U121 ( .A(n95), .B(n100), .C(ena[2]), .D(q[8]), .E(q[11]), .Z(
        n91) );
  GTECH_NOT U122 ( .A(q[9]), .Z(n100) );
  GTECH_NOT U123 ( .A(q[10]), .Z(n95) );
  GTECH_NOT U124 ( .A(n105), .Z(ena[2]) );
  GTECH_MUX2 U125 ( .A(n106), .B(n107), .S(q[7]), .Z(N26) );
  GTECH_AO21 U126 ( .A(n108), .B(n109), .C(n110), .Z(n107) );
  GTECH_AND2 U127 ( .A(q[6]), .B(n111), .Z(n106) );
  GTECH_NAND3 U128 ( .A(n105), .B(n89), .C(n112), .Z(N25) );
  GTECH_MUX2 U129 ( .A(n111), .B(n110), .S(q[6]), .Z(N24) );
  GTECH_AO21 U130 ( .A(n108), .B(n113), .C(N22), .Z(n110) );
  GTECH_NOT U131 ( .A(n114), .Z(n111) );
  GTECH_NAND3 U132 ( .A(n108), .B(q[4]), .C(q[5]), .Z(n114) );
  GTECH_MUX2 U133 ( .A(n115), .B(N22), .S(q[5]), .Z(N23) );
  GTECH_AND2 U134 ( .A(n108), .B(q[4]), .Z(n115) );
  GTECH_NOT U135 ( .A(n116), .Z(N22) );
  GTECH_NAND2 U136 ( .A(n108), .B(n117), .Z(n116) );
  GTECH_NOT U137 ( .A(q[4]), .Z(n117) );
  GTECH_NOT U138 ( .A(n112), .Z(n108) );
  GTECH_NAND3 U139 ( .A(n105), .B(n89), .C(ena[1]), .Z(n112) );
  GTECH_NAND5 U140 ( .A(n113), .B(n109), .C(ena[1]), .D(q[7]), .E(q[4]), .Z(
        n105) );
  GTECH_NOT U141 ( .A(n118), .Z(ena[1]) );
  GTECH_NOT U142 ( .A(q[6]), .Z(n109) );
  GTECH_NOT U143 ( .A(q[5]), .Z(n113) );
  GTECH_MUX2 U144 ( .A(n119), .B(n120), .S(q[3]), .Z(N13) );
  GTECH_AO21 U145 ( .A(n121), .B(n122), .C(n123), .Z(n120) );
  GTECH_AND2 U146 ( .A(q[2]), .B(n124), .Z(n119) );
  GTECH_MUX2 U147 ( .A(n124), .B(n123), .S(q[2]), .Z(N12) );
  GTECH_AO21 U148 ( .A(n121), .B(n125), .C(N10), .Z(n123) );
  GTECH_NOT U149 ( .A(n126), .Z(n124) );
  GTECH_NAND3 U150 ( .A(n121), .B(q[0]), .C(q[1]), .Z(n126) );
  GTECH_MUX2 U151 ( .A(n127), .B(N10), .S(q[1]), .Z(N11) );
  GTECH_AND2 U152 ( .A(n121), .B(q[0]), .Z(n127) );
  GTECH_NOT U153 ( .A(n128), .Z(N10) );
  GTECH_NAND2 U154 ( .A(n121), .B(n129), .Z(n128) );
  GTECH_NOT U155 ( .A(q[0]), .Z(n129) );
  GTECH_NOT U156 ( .A(n130), .Z(n121) );
  GTECH_NAND2 U157 ( .A(n118), .B(n89), .Z(n130) );
  GTECH_NOT U158 ( .A(reset), .Z(n89) );
  GTECH_NAND4 U159 ( .A(q[3]), .B(q[0]), .C(n125), .D(n122), .Z(n118) );
  GTECH_NOT U160 ( .A(q[2]), .Z(n122) );
  GTECH_NOT U161 ( .A(q[1]), .Z(n125) );
endmodule

