
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127;

  GTECH_XOR2 U82 ( .A(n63), .B(n64), .Z(sum[9]) );
  GTECH_XOR2 U83 ( .A(n65), .B(n66), .Z(sum[8]) );
  GTECH_XNOR2 U84 ( .A(n67), .B(n68), .Z(sum[7]) );
  GTECH_AOI21 U85 ( .A(n69), .B(n70), .C(n71), .Z(n68) );
  GTECH_XOR2 U86 ( .A(n70), .B(n69), .Z(sum[6]) );
  GTECH_AO22 U87 ( .A(b[5]), .B(a[5]), .C(n72), .D(n73), .Z(n69) );
  GTECH_XOR2 U88 ( .A(n73), .B(n72), .Z(sum[5]) );
  GTECH_AO22 U89 ( .A(n74), .B(n75), .C(b[4]), .D(a[4]), .Z(n72) );
  GTECH_XOR2 U90 ( .A(n75), .B(n74), .Z(sum[4]) );
  GTECH_XNOR2 U91 ( .A(n76), .B(n77), .Z(sum[3]) );
  GTECH_AOI21 U92 ( .A(n78), .B(n79), .C(n80), .Z(n77) );
  GTECH_XNOR2 U93 ( .A(n81), .B(n78), .Z(sum[2]) );
  GTECH_AO21 U94 ( .A(n82), .B(n83), .C(n84), .Z(n78) );
  GTECH_NOT U95 ( .A(n85), .Z(n84) );
  GTECH_XOR2 U96 ( .A(n82), .B(n83), .Z(sum[1]) );
  GTECH_AO22 U97 ( .A(n86), .B(cin), .C(a[0]), .D(b[0]), .Z(n83) );
  GTECH_XNOR2 U98 ( .A(n87), .B(n88), .Z(sum[15]) );
  GTECH_AOI21 U99 ( .A(n89), .B(n90), .C(n91), .Z(n88) );
  GTECH_XOR2 U100 ( .A(n90), .B(n89), .Z(sum[14]) );
  GTECH_AO22 U101 ( .A(n92), .B(n93), .C(b[13]), .D(a[13]), .Z(n89) );
  GTECH_XOR2 U102 ( .A(n93), .B(n92), .Z(sum[13]) );
  GTECH_AO22 U103 ( .A(a[12]), .B(b[12]), .C(cout), .D(n94), .Z(n92) );
  GTECH_XOR2 U104 ( .A(n94), .B(cout), .Z(sum[12]) );
  GTECH_XOR2 U105 ( .A(n95), .B(n96), .Z(sum[11]) );
  GTECH_OA21 U106 ( .A(n97), .B(n98), .C(n99), .Z(n96) );
  GTECH_XNOR2 U107 ( .A(n100), .B(n97), .Z(sum[10]) );
  GTECH_AOI21 U108 ( .A(n63), .B(n64), .C(n101), .Z(n97) );
  GTECH_AO21 U109 ( .A(n65), .B(n66), .C(n102), .Z(n64) );
  GTECH_XOR2 U110 ( .A(cin), .B(n86), .Z(sum[0]) );
  GTECH_AO21 U111 ( .A(n103), .B(n66), .C(n104), .Z(cout) );
  GTECH_AO21 U112 ( .A(n105), .B(n74), .C(n106), .Z(n66) );
  GTECH_AO21 U113 ( .A(cin), .B(n107), .C(n108), .Z(n74) );
  GTECH_AND3 U114 ( .A(n105), .B(n107), .C(n103), .Z(Pm) );
  GTECH_NOT U115 ( .A(n109), .Z(n107) );
  GTECH_NAND5 U116 ( .A(n79), .B(n82), .C(n76), .D(n110), .E(n86), .Z(n109) );
  GTECH_XOR2 U117 ( .A(a[0]), .B(b[0]), .Z(n86) );
  GTECH_AO21 U118 ( .A(n103), .B(n111), .C(n104), .Z(Gm) );
  GTECH_AO22 U119 ( .A(b[15]), .B(a[15]), .C(n112), .D(n87), .Z(n104) );
  GTECH_AO21 U120 ( .A(n113), .B(n90), .C(n91), .Z(n112) );
  GTECH_AND2 U121 ( .A(a[14]), .B(b[14]), .Z(n91) );
  GTECH_AO21 U122 ( .A(b[13]), .B(a[13]), .C(n114), .Z(n113) );
  GTECH_AND3 U123 ( .A(a[12]), .B(n93), .C(b[12]), .Z(n114) );
  GTECH_AO21 U124 ( .A(n105), .B(n108), .C(n106), .Z(n111) );
  GTECH_OAI2N2 U125 ( .A(n115), .B(n95), .C(b[11]), .D(a[11]), .Z(n106) );
  GTECH_OA21 U126 ( .A(n116), .B(n98), .C(n99), .Z(n115) );
  GTECH_AOI21 U127 ( .A(n63), .B(n102), .C(n101), .Z(n116) );
  GTECH_AND2 U128 ( .A(a[9]), .B(b[9]), .Z(n101) );
  GTECH_NOT U129 ( .A(n117), .Z(n108) );
  GTECH_AOI222 U130 ( .A(a[7]), .B(b[7]), .C(n110), .D(n118), .E(n67), .F(n119), .Z(n117) );
  GTECH_AO21 U131 ( .A(n70), .B(n120), .C(n71), .Z(n119) );
  GTECH_AND2 U132 ( .A(b[6]), .B(a[6]), .Z(n71) );
  GTECH_AO22 U133 ( .A(a[4]), .B(n121), .C(b[5]), .D(a[5]), .Z(n120) );
  GTECH_AND2 U134 ( .A(n73), .B(b[4]), .Z(n121) );
  GTECH_AO22 U135 ( .A(n122), .B(n76), .C(b[3]), .D(a[3]), .Z(n118) );
  GTECH_XOR2 U136 ( .A(a[3]), .B(b[3]), .Z(n76) );
  GTECH_OR_NOT U137 ( .A(n80), .B(n123), .Z(n122) );
  GTECH_AO21 U138 ( .A(n85), .B(n124), .C(n81), .Z(n123) );
  GTECH_NOT U139 ( .A(n79), .Z(n81) );
  GTECH_XOR2 U140 ( .A(a[2]), .B(b[2]), .Z(n79) );
  GTECH_NAND3 U141 ( .A(a[0]), .B(n82), .C(b[0]), .Z(n124) );
  GTECH_XOR2 U142 ( .A(a[1]), .B(b[1]), .Z(n82) );
  GTECH_NAND2 U143 ( .A(a[1]), .B(b[1]), .Z(n85) );
  GTECH_AND2 U144 ( .A(a[2]), .B(b[2]), .Z(n80) );
  GTECH_AND4 U145 ( .A(n75), .B(n73), .C(n70), .D(n67), .Z(n110) );
  GTECH_XOR2 U146 ( .A(a[7]), .B(b[7]), .Z(n67) );
  GTECH_XOR2 U147 ( .A(a[6]), .B(b[6]), .Z(n70) );
  GTECH_XOR2 U148 ( .A(a[5]), .B(b[5]), .Z(n73) );
  GTECH_XOR2 U149 ( .A(a[4]), .B(b[4]), .Z(n75) );
  GTECH_NOR4 U150 ( .A(n125), .B(n98), .C(n95), .D(n126), .Z(n105) );
  GTECH_NOT U151 ( .A(n63), .Z(n126) );
  GTECH_XOR2 U152 ( .A(a[9]), .B(b[9]), .Z(n63) );
  GTECH_XNOR2 U153 ( .A(a[11]), .B(b[11]), .Z(n95) );
  GTECH_NOT U154 ( .A(n100), .Z(n98) );
  GTECH_OA21 U155 ( .A(a[10]), .B(b[10]), .C(n99), .Z(n100) );
  GTECH_NAND2 U156 ( .A(b[10]), .B(a[10]), .Z(n99) );
  GTECH_NOT U157 ( .A(n65), .Z(n125) );
  GTECH_OA21 U158 ( .A(a[8]), .B(b[8]), .C(n127), .Z(n65) );
  GTECH_NOT U159 ( .A(n102), .Z(n127) );
  GTECH_AND2 U160 ( .A(b[8]), .B(a[8]), .Z(n102) );
  GTECH_AND4 U161 ( .A(n94), .B(n87), .C(n90), .D(n93), .Z(n103) );
  GTECH_XOR2 U162 ( .A(a[13]), .B(b[13]), .Z(n93) );
  GTECH_XOR2 U163 ( .A(a[14]), .B(b[14]), .Z(n90) );
  GTECH_XOR2 U164 ( .A(a[15]), .B(b[15]), .Z(n87) );
  GTECH_XOR2 U165 ( .A(a[12]), .B(b[12]), .Z(n94) );
endmodule

