
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144;

  GTECH_XOR2 U89 ( .A(n70), .B(n71), .Z(sum[9]) );
  GTECH_XNOR2 U90 ( .A(n72), .B(n73), .Z(sum[8]) );
  GTECH_XNOR2 U91 ( .A(n74), .B(n75), .Z(sum[7]) );
  GTECH_OA21 U92 ( .A(n76), .B(n77), .C(n78), .Z(n75) );
  GTECH_XNOR2 U93 ( .A(n76), .B(n79), .Z(sum[6]) );
  GTECH_OA21 U94 ( .A(n80), .B(n81), .C(n82), .Z(n76) );
  GTECH_XOR2 U95 ( .A(n81), .B(n80), .Z(sum[5]) );
  GTECH_AOI22 U96 ( .A(b[4]), .B(a[4]), .C(n83), .D(n84), .Z(n80) );
  GTECH_NOT U97 ( .A(n85), .Z(n81) );
  GTECH_XNOR2 U98 ( .A(n84), .B(n86), .Z(sum[4]) );
  GTECH_XNOR2 U99 ( .A(n87), .B(n88), .Z(sum[3]) );
  GTECH_OA21 U100 ( .A(n89), .B(n90), .C(n91), .Z(n88) );
  GTECH_XNOR2 U101 ( .A(n92), .B(n89), .Z(sum[2]) );
  GTECH_AOI21 U102 ( .A(n93), .B(n94), .C(n95), .Z(n89) );
  GTECH_XOR2 U103 ( .A(n94), .B(n93), .Z(sum[1]) );
  GTECH_NOT U104 ( .A(n96), .Z(n93) );
  GTECH_AOI21 U105 ( .A(n97), .B(cin), .C(n98), .Z(n96) );
  GTECH_XNOR2 U106 ( .A(n99), .B(n100), .Z(sum[15]) );
  GTECH_AOI21 U107 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_XOR2 U108 ( .A(n101), .B(n102), .Z(sum[14]) );
  GTECH_NOT U109 ( .A(n104), .Z(n101) );
  GTECH_AOI21 U110 ( .A(n105), .B(n106), .C(n107), .Z(n104) );
  GTECH_XOR2 U111 ( .A(n106), .B(n105), .Z(sum[13]) );
  GTECH_AO22 U112 ( .A(cout), .B(n108), .C(a[12]), .D(b[12]), .Z(n105) );
  GTECH_XNOR2 U113 ( .A(n108), .B(n109), .Z(sum[12]) );
  GTECH_XOR2 U114 ( .A(n110), .B(n111), .Z(sum[11]) );
  GTECH_OA21 U115 ( .A(n112), .B(n113), .C(n114), .Z(n111) );
  GTECH_XOR2 U116 ( .A(n112), .B(n113), .Z(sum[10]) );
  GTECH_OA21 U117 ( .A(n71), .B(n70), .C(n115), .Z(n112) );
  GTECH_OA21 U118 ( .A(n73), .B(n116), .C(n117), .Z(n71) );
  GTECH_XOR2 U119 ( .A(cin), .B(n97), .Z(sum[0]) );
  GTECH_NOT U120 ( .A(n109), .Z(cout) );
  GTECH_OA21 U121 ( .A(n73), .B(n118), .C(n119), .Z(n109) );
  GTECH_AOI21 U122 ( .A(n83), .B(n120), .C(n121), .Z(n73) );
  GTECH_NOT U123 ( .A(n86), .Z(n83) );
  GTECH_AOI21 U124 ( .A(n122), .B(cin), .C(n123), .Z(n86) );
  GTECH_AND3 U125 ( .A(n120), .B(n122), .C(n124), .Z(Pm) );
  GTECH_AND5 U126 ( .A(n87), .B(n94), .C(n97), .D(n125), .E(n92), .Z(n122) );
  GTECH_XOR2 U127 ( .A(a[0]), .B(b[0]), .Z(n97) );
  GTECH_NOT U128 ( .A(n126), .Z(Gm) );
  GTECH_OA21 U129 ( .A(n127), .B(n118), .C(n119), .Z(n126) );
  GTECH_AND_NOT U130 ( .A(n128), .B(n129), .Z(n119) );
  GTECH_OA21 U131 ( .A(n103), .B(n130), .C(n99), .Z(n129) );
  GTECH_OA21 U132 ( .A(n131), .B(n107), .C(n102), .Z(n130) );
  GTECH_AND2 U133 ( .A(a[13]), .B(b[13]), .Z(n107) );
  GTECH_AND3 U134 ( .A(a[12]), .B(n106), .C(b[12]), .Z(n131) );
  GTECH_NOT U135 ( .A(n124), .Z(n118) );
  GTECH_AND4 U136 ( .A(n99), .B(n102), .C(n108), .D(n106), .Z(n124) );
  GTECH_XOR2 U137 ( .A(a[13]), .B(b[13]), .Z(n106) );
  GTECH_XOR2 U138 ( .A(a[12]), .B(b[12]), .Z(n108) );
  GTECH_OA21 U139 ( .A(a[14]), .B(b[14]), .C(n132), .Z(n102) );
  GTECH_NOT U140 ( .A(n103), .Z(n132) );
  GTECH_AND2 U141 ( .A(a[14]), .B(b[14]), .Z(n103) );
  GTECH_OA21 U142 ( .A(b[15]), .B(a[15]), .C(n128), .Z(n99) );
  GTECH_NAND2 U143 ( .A(a[15]), .B(b[15]), .Z(n128) );
  GTECH_AOI21 U144 ( .A(n123), .B(n120), .C(n121), .Z(n127) );
  GTECH_OAI2N2 U145 ( .A(n133), .B(n110), .C(b[11]), .D(a[11]), .Z(n121) );
  GTECH_OA21 U146 ( .A(n134), .B(n113), .C(n114), .Z(n133) );
  GTECH_OA21 U147 ( .A(n70), .B(n117), .C(n115), .Z(n134) );
  GTECH_NAND2 U148 ( .A(b[9]), .B(a[9]), .Z(n115) );
  GTECH_NOR4 U149 ( .A(n116), .B(n113), .C(n110), .D(n70), .Z(n120) );
  GTECH_XNOR2 U150 ( .A(a[9]), .B(b[9]), .Z(n70) );
  GTECH_XNOR2 U151 ( .A(a[11]), .B(b[11]), .Z(n110) );
  GTECH_NOT U152 ( .A(n135), .Z(n113) );
  GTECH_OA21 U153 ( .A(a[10]), .B(b[10]), .C(n114), .Z(n135) );
  GTECH_NAND2 U154 ( .A(a[10]), .B(b[10]), .Z(n114) );
  GTECH_NOT U155 ( .A(n72), .Z(n116) );
  GTECH_OA21 U156 ( .A(b[8]), .B(a[8]), .C(n117), .Z(n72) );
  GTECH_NAND2 U157 ( .A(a[8]), .B(b[8]), .Z(n117) );
  GTECH_NOT U158 ( .A(n136), .Z(n123) );
  GTECH_AOI222 U159 ( .A(a[7]), .B(b[7]), .C(n125), .D(n137), .E(n74), .F(n138), .Z(n136) );
  GTECH_OR_NOT U160 ( .A(n139), .B(n78), .Z(n138) );
  GTECH_AOI21 U161 ( .A(n140), .B(n82), .C(n77), .Z(n139) );
  GTECH_NOT U162 ( .A(n79), .Z(n77) );
  GTECH_NAND2 U163 ( .A(b[5]), .B(a[5]), .Z(n82) );
  GTECH_NAND3 U164 ( .A(b[4]), .B(n85), .C(a[4]), .Z(n140) );
  GTECH_OAI2N2 U165 ( .A(n141), .B(n142), .C(b[3]), .D(a[3]), .Z(n137) );
  GTECH_NOT U166 ( .A(n87), .Z(n142) );
  GTECH_XOR2 U167 ( .A(a[3]), .B(b[3]), .Z(n87) );
  GTECH_OA21 U168 ( .A(n143), .B(n90), .C(n91), .Z(n141) );
  GTECH_NOT U169 ( .A(n92), .Z(n90) );
  GTECH_OA21 U170 ( .A(b[2]), .B(a[2]), .C(n91), .Z(n92) );
  GTECH_NAND2 U171 ( .A(a[2]), .B(b[2]), .Z(n91) );
  GTECH_AOI21 U172 ( .A(n94), .B(n98), .C(n95), .Z(n143) );
  GTECH_NOT U173 ( .A(n144), .Z(n95) );
  GTECH_NAND2 U174 ( .A(a[1]), .B(b[1]), .Z(n144) );
  GTECH_AND2 U175 ( .A(a[0]), .B(b[0]), .Z(n98) );
  GTECH_XOR2 U176 ( .A(a[1]), .B(b[1]), .Z(n94) );
  GTECH_AND4 U177 ( .A(n79), .B(n84), .C(n74), .D(n85), .Z(n125) );
  GTECH_XOR2 U178 ( .A(a[5]), .B(b[5]), .Z(n85) );
  GTECH_XOR2 U179 ( .A(a[7]), .B(b[7]), .Z(n74) );
  GTECH_XOR2 U180 ( .A(a[4]), .B(b[4]), .Z(n84) );
  GTECH_OA21 U181 ( .A(a[6]), .B(b[6]), .C(n78), .Z(n79) );
  GTECH_NAND2 U182 ( .A(a[6]), .B(b[6]), .Z(n78) );
endmodule

