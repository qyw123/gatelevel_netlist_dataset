
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n85) );
  GTECH_XNOR2 U78 ( .A(n84), .B(n90), .Z(N154) );
  GTECH_XNOR2 U79 ( .A(n91), .B(n92), .Z(n90) );
  GTECH_NOT U80 ( .A(n86), .Z(n92) );
  GTECH_XNOR2 U81 ( .A(n93), .B(n88), .Z(n86) );
  GTECH_NOT U82 ( .A(n94), .Z(n88) );
  GTECH_NAND2 U83 ( .A(I_b[7]), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U84 ( .A(n89), .Z(n93) );
  GTECH_OAI21 U85 ( .A(n95), .B(n96), .C(n97), .Z(n89) );
  GTECH_OAI21 U86 ( .A(n98), .B(n99), .C(n100), .Z(n97) );
  GTECH_NOT U87 ( .A(n99), .Z(n95) );
  GTECH_NOT U88 ( .A(n87), .Z(n91) );
  GTECH_OAI2N2 U89 ( .A(n101), .B(n102), .C(n103), .D(n104), .Z(n87) );
  GTECH_NAND2 U90 ( .A(n101), .B(n102), .Z(n104) );
  GTECH_NOT U91 ( .A(n105), .Z(n84) );
  GTECH_NAND2 U92 ( .A(n106), .B(n107), .Z(n105) );
  GTECH_NOT U93 ( .A(n108), .Z(n106) );
  GTECH_XNOR2 U94 ( .A(n107), .B(n108), .Z(N153) );
  GTECH_XOR3 U95 ( .A(n109), .B(n101), .C(n103), .Z(n108) );
  GTECH_XOR3 U96 ( .A(n98), .B(n100), .C(n99), .Z(n103) );
  GTECH_OAI21 U97 ( .A(n110), .B(n111), .C(n112), .Z(n99) );
  GTECH_OAI21 U98 ( .A(n113), .B(n114), .C(n115), .Z(n112) );
  GTECH_NOT U99 ( .A(n114), .Z(n110) );
  GTECH_NOT U100 ( .A(n116), .Z(n100) );
  GTECH_NAND2 U101 ( .A(I_b[7]), .B(I_a[6]), .Z(n116) );
  GTECH_NOT U102 ( .A(n96), .Z(n98) );
  GTECH_NAND2 U103 ( .A(I_a[7]), .B(I_b[6]), .Z(n96) );
  GTECH_ADD_ABC U104 ( .A(n117), .B(n118), .C(n119), .COUT(n101) );
  GTECH_NOT U105 ( .A(n120), .Z(n119) );
  GTECH_XNOR2 U106 ( .A(n121), .B(n122), .Z(n118) );
  GTECH_NAND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n122) );
  GTECH_NOT U108 ( .A(n102), .Z(n109) );
  GTECH_NAND2 U109 ( .A(I_a[7]), .B(n123), .Z(n102) );
  GTECH_NOT U110 ( .A(n124), .Z(n107) );
  GTECH_NAND2 U111 ( .A(n125), .B(n126), .Z(n124) );
  GTECH_NOT U112 ( .A(n127), .Z(n126) );
  GTECH_XNOR2 U113 ( .A(n127), .B(n125), .Z(N152) );
  GTECH_XOR4 U114 ( .A(n121), .B(n128), .C(n117), .D(n120), .Z(n125) );
  GTECH_XOR3 U115 ( .A(n113), .B(n115), .C(n114), .Z(n120) );
  GTECH_OAI21 U116 ( .A(n129), .B(n130), .C(n131), .Z(n114) );
  GTECH_OAI21 U117 ( .A(n132), .B(n133), .C(n134), .Z(n131) );
  GTECH_NOT U118 ( .A(n133), .Z(n129) );
  GTECH_NOT U119 ( .A(n135), .Z(n115) );
  GTECH_NAND2 U120 ( .A(I_b[7]), .B(I_a[5]), .Z(n135) );
  GTECH_NOT U121 ( .A(n111), .Z(n113) );
  GTECH_NAND2 U122 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_ADD_ABC U123 ( .A(n136), .B(n137), .C(n138), .COUT(n117) );
  GTECH_NOT U124 ( .A(n139), .Z(n138) );
  GTECH_XOR3 U125 ( .A(n140), .B(n141), .C(n142), .Z(n137) );
  GTECH_AND2 U126 ( .A(I_a[7]), .B(I_b[5]), .Z(n128) );
  GTECH_NOT U127 ( .A(n123), .Z(n121) );
  GTECH_OAI21 U128 ( .A(n142), .B(n143), .C(n144), .Z(n123) );
  GTECH_OAI21 U129 ( .A(n140), .B(n145), .C(n141), .Z(n144) );
  GTECH_NOT U130 ( .A(n143), .Z(n140) );
  GTECH_NOT U131 ( .A(n145), .Z(n142) );
  GTECH_ADD_ABC U132 ( .A(n146), .B(n147), .C(n148), .COUT(n127) );
  GTECH_NOT U133 ( .A(n149), .Z(n148) );
  GTECH_AOI2N2 U134 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n147) );
  GTECH_OA21 U135 ( .A(n154), .B(n155), .C(n156), .Z(n146) );
  GTECH_XOR3 U136 ( .A(n157), .B(n149), .C(n158), .Z(N151) );
  GTECH_OA21 U137 ( .A(n154), .B(n155), .C(n156), .Z(n158) );
  GTECH_OAI21 U138 ( .A(n159), .B(n160), .C(n161), .Z(n156) );
  GTECH_XOR3 U139 ( .A(n139), .B(n136), .C(n162), .Z(n149) );
  GTECH_XOR3 U140 ( .A(n141), .B(n145), .C(n143), .Z(n162) );
  GTECH_NAND2 U141 ( .A(I_a[7]), .B(I_b[4]), .Z(n143) );
  GTECH_OAI21 U142 ( .A(n163), .B(n164), .C(n165), .Z(n145) );
  GTECH_OAI21 U143 ( .A(n166), .B(n167), .C(n168), .Z(n165) );
  GTECH_NOT U144 ( .A(n169), .Z(n141) );
  GTECH_NAND2 U145 ( .A(I_a[6]), .B(I_b[5]), .Z(n169) );
  GTECH_ADD_ABC U146 ( .A(n170), .B(n171), .C(n172), .COUT(n136) );
  GTECH_NOT U147 ( .A(n173), .Z(n172) );
  GTECH_XOR3 U148 ( .A(n166), .B(n168), .C(n163), .Z(n171) );
  GTECH_NOT U149 ( .A(n167), .Z(n163) );
  GTECH_NOT U150 ( .A(n164), .Z(n166) );
  GTECH_XOR3 U151 ( .A(n132), .B(n134), .C(n133), .Z(n139) );
  GTECH_OAI21 U152 ( .A(n174), .B(n175), .C(n176), .Z(n133) );
  GTECH_OAI21 U153 ( .A(n177), .B(n178), .C(n179), .Z(n176) );
  GTECH_NOT U154 ( .A(n178), .Z(n174) );
  GTECH_NOT U155 ( .A(n180), .Z(n134) );
  GTECH_NAND2 U156 ( .A(I_b[7]), .B(I_a[4]), .Z(n180) );
  GTECH_NOT U157 ( .A(n130), .Z(n132) );
  GTECH_NAND2 U158 ( .A(I_b[6]), .B(I_a[5]), .Z(n130) );
  GTECH_AOI2N2 U159 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n157) );
  GTECH_NOT U160 ( .A(I_a[7]), .Z(n153) );
  GTECH_XOR3 U161 ( .A(n154), .B(n159), .C(n181), .Z(N150) );
  GTECH_NOT U162 ( .A(n161), .Z(n181) );
  GTECH_XOR3 U163 ( .A(n173), .B(n170), .C(n182), .Z(n161) );
  GTECH_XOR3 U164 ( .A(n168), .B(n167), .C(n164), .Z(n182) );
  GTECH_NAND2 U165 ( .A(I_a[6]), .B(I_b[4]), .Z(n164) );
  GTECH_OAI21 U166 ( .A(n183), .B(n184), .C(n185), .Z(n167) );
  GTECH_OAI21 U167 ( .A(n186), .B(n187), .C(n188), .Z(n185) );
  GTECH_NOT U168 ( .A(n189), .Z(n168) );
  GTECH_NAND2 U169 ( .A(I_a[5]), .B(I_b[5]), .Z(n189) );
  GTECH_ADD_ABC U170 ( .A(n190), .B(n191), .C(n192), .COUT(n170) );
  GTECH_NOT U171 ( .A(n193), .Z(n192) );
  GTECH_XOR3 U172 ( .A(n186), .B(n188), .C(n183), .Z(n191) );
  GTECH_NOT U173 ( .A(n187), .Z(n183) );
  GTECH_NOT U174 ( .A(n184), .Z(n186) );
  GTECH_XOR3 U175 ( .A(n177), .B(n179), .C(n178), .Z(n173) );
  GTECH_OAI21 U176 ( .A(n194), .B(n195), .C(n196), .Z(n178) );
  GTECH_OAI21 U177 ( .A(n197), .B(n198), .C(n199), .Z(n196) );
  GTECH_NOT U178 ( .A(n198), .Z(n194) );
  GTECH_NOT U179 ( .A(n200), .Z(n179) );
  GTECH_NAND2 U180 ( .A(I_b[7]), .B(I_a[3]), .Z(n200) );
  GTECH_NOT U181 ( .A(n175), .Z(n177) );
  GTECH_NAND2 U182 ( .A(I_b[6]), .B(I_a[4]), .Z(n175) );
  GTECH_NOT U183 ( .A(n155), .Z(n159) );
  GTECH_XNOR2 U184 ( .A(n201), .B(n202), .Z(n155) );
  GTECH_NOT U185 ( .A(n150), .Z(n202) );
  GTECH_XNOR2 U186 ( .A(n152), .B(n203), .Z(n150) );
  GTECH_AND2 U187 ( .A(I_a[7]), .B(I_b[3]), .Z(n203) );
  GTECH_AND2 U188 ( .A(n204), .B(n205), .Z(n152) );
  GTECH_OR_NOT U189 ( .A(n206), .B(n207), .Z(n205) );
  GTECH_OAI21 U190 ( .A(n208), .B(n207), .C(n209), .Z(n204) );
  GTECH_NOT U191 ( .A(n151), .Z(n201) );
  GTECH_OAI2N2 U192 ( .A(n210), .B(n211), .C(n212), .D(n213), .Z(n151) );
  GTECH_NAND2 U193 ( .A(n210), .B(n211), .Z(n213) );
  GTECH_NOT U194 ( .A(n160), .Z(n154) );
  GTECH_OAI2N2 U195 ( .A(n214), .B(n215), .C(n216), .D(n217), .Z(n160) );
  GTECH_NAND2 U196 ( .A(n214), .B(n215), .Z(n217) );
  GTECH_XOR3 U197 ( .A(n214), .B(n218), .C(n219), .Z(N149) );
  GTECH_NOT U198 ( .A(n216), .Z(n219) );
  GTECH_XOR3 U199 ( .A(n193), .B(n190), .C(n220), .Z(n216) );
  GTECH_XOR3 U200 ( .A(n188), .B(n187), .C(n184), .Z(n220) );
  GTECH_NAND2 U201 ( .A(I_a[5]), .B(I_b[4]), .Z(n184) );
  GTECH_OAI21 U202 ( .A(n221), .B(n222), .C(n223), .Z(n187) );
  GTECH_OAI21 U203 ( .A(n224), .B(n225), .C(n226), .Z(n223) );
  GTECH_NOT U204 ( .A(n227), .Z(n188) );
  GTECH_NAND2 U205 ( .A(I_b[5]), .B(I_a[4]), .Z(n227) );
  GTECH_ADD_ABC U206 ( .A(n228), .B(n229), .C(n230), .COUT(n190) );
  GTECH_XOR3 U207 ( .A(n224), .B(n226), .C(n221), .Z(n229) );
  GTECH_NOT U208 ( .A(n225), .Z(n221) );
  GTECH_OA21 U209 ( .A(n231), .B(n232), .C(n233), .Z(n228) );
  GTECH_XOR3 U210 ( .A(n197), .B(n199), .C(n198), .Z(n193) );
  GTECH_OAI21 U211 ( .A(n234), .B(n235), .C(n236), .Z(n198) );
  GTECH_NOT U212 ( .A(n237), .Z(n199) );
  GTECH_NAND2 U213 ( .A(I_b[7]), .B(I_a[2]), .Z(n237) );
  GTECH_NOT U214 ( .A(n195), .Z(n197) );
  GTECH_NAND2 U215 ( .A(I_b[6]), .B(I_a[3]), .Z(n195) );
  GTECH_NOT U216 ( .A(n215), .Z(n218) );
  GTECH_XOR3 U217 ( .A(n238), .B(n210), .C(n212), .Z(n215) );
  GTECH_XOR3 U218 ( .A(n208), .B(n209), .C(n207), .Z(n212) );
  GTECH_OAI21 U219 ( .A(n239), .B(n240), .C(n241), .Z(n207) );
  GTECH_OAI21 U220 ( .A(n242), .B(n243), .C(n244), .Z(n241) );
  GTECH_NOT U221 ( .A(n243), .Z(n239) );
  GTECH_NOT U222 ( .A(n245), .Z(n209) );
  GTECH_NAND2 U223 ( .A(I_a[6]), .B(I_b[3]), .Z(n245) );
  GTECH_NOT U224 ( .A(n206), .Z(n208) );
  GTECH_NAND2 U225 ( .A(I_a[7]), .B(I_b[2]), .Z(n206) );
  GTECH_ADD_ABC U226 ( .A(n246), .B(n247), .C(n248), .COUT(n210) );
  GTECH_XNOR2 U227 ( .A(n249), .B(n250), .Z(n247) );
  GTECH_NAND2 U228 ( .A(I_a[7]), .B(I_b[1]), .Z(n250) );
  GTECH_NOT U229 ( .A(n211), .Z(n238) );
  GTECH_NAND2 U230 ( .A(I_a[7]), .B(n251), .Z(n211) );
  GTECH_ADD_ABC U231 ( .A(n252), .B(n253), .C(n254), .COUT(n214) );
  GTECH_XOR3 U232 ( .A(n246), .B(n255), .C(n248), .Z(n253) );
  GTECH_NOT U233 ( .A(n256), .Z(n248) );
  GTECH_XOR3 U234 ( .A(n257), .B(n254), .C(n252), .Z(N148) );
  GTECH_ADD_ABC U235 ( .A(n258), .B(n259), .C(n260), .COUT(n252) );
  GTECH_NOT U236 ( .A(n261), .Z(n260) );
  GTECH_XOR3 U237 ( .A(n262), .B(n263), .C(n264), .Z(n259) );
  GTECH_NOT U238 ( .A(n265), .Z(n263) );
  GTECH_XOR3 U239 ( .A(n266), .B(n230), .C(n267), .Z(n254) );
  GTECH_OAI21 U240 ( .A(n231), .B(n232), .C(n233), .Z(n267) );
  GTECH_OAI21 U241 ( .A(n268), .B(n269), .C(n270), .Z(n233) );
  GTECH_NOT U242 ( .A(n231), .Z(n269) );
  GTECH_XOR3 U243 ( .A(n271), .B(n272), .C(n236), .Z(n230) );
  GTECH_NAND3 U244 ( .A(I_b[6]), .B(I_a[1]), .C(n273), .Z(n236) );
  GTECH_NOT U245 ( .A(n235), .Z(n272) );
  GTECH_NAND2 U246 ( .A(I_b[7]), .B(I_a[1]), .Z(n235) );
  GTECH_NOT U247 ( .A(n234), .Z(n271) );
  GTECH_NAND2 U248 ( .A(I_b[6]), .B(I_a[2]), .Z(n234) );
  GTECH_XOR3 U249 ( .A(n226), .B(n225), .C(n224), .Z(n266) );
  GTECH_NOT U250 ( .A(n222), .Z(n224) );
  GTECH_NAND2 U251 ( .A(I_b[4]), .B(I_a[4]), .Z(n222) );
  GTECH_OAI21 U252 ( .A(n274), .B(n275), .C(n276), .Z(n225) );
  GTECH_OAI21 U253 ( .A(n277), .B(n278), .C(n279), .Z(n276) );
  GTECH_NOT U254 ( .A(n278), .Z(n274) );
  GTECH_NOT U255 ( .A(n280), .Z(n226) );
  GTECH_NAND2 U256 ( .A(I_b[5]), .B(I_a[3]), .Z(n280) );
  GTECH_XOR3 U257 ( .A(n255), .B(n256), .C(n246), .Z(n257) );
  GTECH_ADD_ABC U258 ( .A(n262), .B(n281), .C(n264), .COUT(n246) );
  GTECH_NOT U259 ( .A(n282), .Z(n264) );
  GTECH_XOR3 U260 ( .A(n283), .B(n284), .C(n285), .Z(n281) );
  GTECH_XOR3 U261 ( .A(n242), .B(n244), .C(n243), .Z(n256) );
  GTECH_OAI21 U262 ( .A(n286), .B(n287), .C(n288), .Z(n243) );
  GTECH_OAI21 U263 ( .A(n289), .B(n290), .C(n291), .Z(n288) );
  GTECH_NOT U264 ( .A(n290), .Z(n286) );
  GTECH_NOT U265 ( .A(n292), .Z(n244) );
  GTECH_NAND2 U266 ( .A(I_a[5]), .B(I_b[3]), .Z(n292) );
  GTECH_NOT U267 ( .A(n240), .Z(n242) );
  GTECH_NAND2 U268 ( .A(I_a[6]), .B(I_b[2]), .Z(n240) );
  GTECH_XNOR2 U269 ( .A(n249), .B(n293), .Z(n255) );
  GTECH_NAND2 U270 ( .A(I_a[7]), .B(I_b[1]), .Z(n293) );
  GTECH_NOT U271 ( .A(n251), .Z(n249) );
  GTECH_OAI21 U272 ( .A(n285), .B(n294), .C(n295), .Z(n251) );
  GTECH_OAI21 U273 ( .A(n283), .B(n296), .C(n284), .Z(n295) );
  GTECH_NOT U274 ( .A(n296), .Z(n285) );
  GTECH_XOR3 U275 ( .A(n261), .B(n258), .C(n297), .Z(N147) );
  GTECH_XOR3 U276 ( .A(n282), .B(n262), .C(n265), .Z(n297) );
  GTECH_XOR3 U277 ( .A(n283), .B(n284), .C(n296), .Z(n265) );
  GTECH_OAI21 U278 ( .A(n298), .B(n299), .C(n300), .Z(n296) );
  GTECH_OAI21 U279 ( .A(n301), .B(n302), .C(n303), .Z(n300) );
  GTECH_NOT U280 ( .A(n304), .Z(n284) );
  GTECH_NAND2 U281 ( .A(I_a[6]), .B(I_b[1]), .Z(n304) );
  GTECH_NOT U282 ( .A(n294), .Z(n283) );
  GTECH_NAND2 U283 ( .A(I_a[7]), .B(I_b[0]), .Z(n294) );
  GTECH_ADD_ABC U284 ( .A(n305), .B(n306), .C(n307), .COUT(n262) );
  GTECH_XOR3 U285 ( .A(n301), .B(n303), .C(n298), .Z(n306) );
  GTECH_NOT U286 ( .A(n302), .Z(n298) );
  GTECH_XOR3 U287 ( .A(n289), .B(n291), .C(n290), .Z(n282) );
  GTECH_OAI21 U288 ( .A(n308), .B(n309), .C(n310), .Z(n290) );
  GTECH_OAI21 U289 ( .A(n311), .B(n312), .C(n313), .Z(n310) );
  GTECH_NOT U290 ( .A(n312), .Z(n308) );
  GTECH_NOT U291 ( .A(n314), .Z(n291) );
  GTECH_NAND2 U292 ( .A(I_b[3]), .B(I_a[4]), .Z(n314) );
  GTECH_NOT U293 ( .A(n287), .Z(n289) );
  GTECH_NAND2 U294 ( .A(I_a[5]), .B(I_b[2]), .Z(n287) );
  GTECH_ADD_ABC U295 ( .A(n315), .B(n316), .C(n317), .COUT(n258) );
  GTECH_XOR3 U296 ( .A(n305), .B(n318), .C(n307), .Z(n316) );
  GTECH_NOT U297 ( .A(n319), .Z(n307) );
  GTECH_OA21 U298 ( .A(n320), .B(n321), .C(n322), .Z(n315) );
  GTECH_XOR3 U299 ( .A(n270), .B(n232), .C(n231), .Z(n261) );
  GTECH_XNOR2 U300 ( .A(n273), .B(n323), .Z(n231) );
  GTECH_AND2 U301 ( .A(I_b[6]), .B(I_a[1]), .Z(n323) );
  GTECH_NOT U302 ( .A(n324), .Z(n273) );
  GTECH_NAND2 U303 ( .A(I_b[7]), .B(I_a[0]), .Z(n324) );
  GTECH_NOT U304 ( .A(n268), .Z(n232) );
  GTECH_XOR3 U305 ( .A(n277), .B(n279), .C(n278), .Z(n268) );
  GTECH_OAI21 U306 ( .A(n325), .B(n326), .C(n327), .Z(n278) );
  GTECH_NOT U307 ( .A(n328), .Z(n279) );
  GTECH_NAND2 U308 ( .A(I_b[5]), .B(I_a[2]), .Z(n328) );
  GTECH_NOT U309 ( .A(n275), .Z(n277) );
  GTECH_NAND2 U310 ( .A(I_b[4]), .B(I_a[3]), .Z(n275) );
  GTECH_NOT U311 ( .A(n329), .Z(n270) );
  GTECH_NAND3 U312 ( .A(I_a[0]), .B(n330), .C(I_b[6]), .Z(n329) );
  GTECH_XOR3 U313 ( .A(n331), .B(n317), .C(n332), .Z(N146) );
  GTECH_OA21 U314 ( .A(n320), .B(n321), .C(n322), .Z(n332) );
  GTECH_OAI21 U315 ( .A(n333), .B(n334), .C(n335), .Z(n322) );
  GTECH_NOT U316 ( .A(n320), .Z(n334) );
  GTECH_XNOR2 U317 ( .A(n336), .B(n330), .Z(n317) );
  GTECH_NOT U318 ( .A(n337), .Z(n330) );
  GTECH_XOR3 U319 ( .A(n338), .B(n339), .C(n327), .Z(n337) );
  GTECH_NAND3 U320 ( .A(I_b[4]), .B(I_a[1]), .C(n340), .Z(n327) );
  GTECH_NOT U321 ( .A(n326), .Z(n339) );
  GTECH_NAND2 U322 ( .A(I_b[5]), .B(I_a[1]), .Z(n326) );
  GTECH_NOT U323 ( .A(n325), .Z(n338) );
  GTECH_NAND2 U324 ( .A(I_b[4]), .B(I_a[2]), .Z(n325) );
  GTECH_AND2 U325 ( .A(I_b[6]), .B(I_a[0]), .Z(n336) );
  GTECH_XOR3 U326 ( .A(n318), .B(n319), .C(n305), .Z(n331) );
  GTECH_ADD_ABC U327 ( .A(n341), .B(n342), .C(n343), .COUT(n305) );
  GTECH_NOT U328 ( .A(n344), .Z(n343) );
  GTECH_XOR3 U329 ( .A(n345), .B(n346), .C(n347), .Z(n342) );
  GTECH_XOR3 U330 ( .A(n311), .B(n313), .C(n312), .Z(n319) );
  GTECH_OAI21 U331 ( .A(n348), .B(n349), .C(n350), .Z(n312) );
  GTECH_OAI21 U332 ( .A(n351), .B(n352), .C(n353), .Z(n350) );
  GTECH_NOT U333 ( .A(n352), .Z(n348) );
  GTECH_NOT U334 ( .A(n354), .Z(n313) );
  GTECH_NAND2 U335 ( .A(I_b[3]), .B(I_a[3]), .Z(n354) );
  GTECH_NOT U336 ( .A(n309), .Z(n311) );
  GTECH_NAND2 U337 ( .A(I_b[2]), .B(I_a[4]), .Z(n309) );
  GTECH_NOT U338 ( .A(n355), .Z(n318) );
  GTECH_XOR3 U339 ( .A(n301), .B(n303), .C(n302), .Z(n355) );
  GTECH_OAI21 U340 ( .A(n347), .B(n356), .C(n357), .Z(n302) );
  GTECH_OAI21 U341 ( .A(n345), .B(n358), .C(n346), .Z(n357) );
  GTECH_NOT U342 ( .A(n356), .Z(n345) );
  GTECH_NOT U343 ( .A(n358), .Z(n347) );
  GTECH_NOT U344 ( .A(n359), .Z(n303) );
  GTECH_NAND2 U345 ( .A(I_a[5]), .B(I_b[1]), .Z(n359) );
  GTECH_NOT U346 ( .A(n299), .Z(n301) );
  GTECH_NAND2 U347 ( .A(I_a[6]), .B(I_b[0]), .Z(n299) );
  GTECH_XOR3 U348 ( .A(n335), .B(n321), .C(n320), .Z(N145) );
  GTECH_XNOR2 U349 ( .A(n340), .B(n360), .Z(n320) );
  GTECH_AND2 U350 ( .A(I_b[4]), .B(I_a[1]), .Z(n360) );
  GTECH_NOT U351 ( .A(n361), .Z(n340) );
  GTECH_NAND2 U352 ( .A(I_b[5]), .B(I_a[0]), .Z(n361) );
  GTECH_NOT U353 ( .A(n333), .Z(n321) );
  GTECH_XOR3 U354 ( .A(n344), .B(n341), .C(n362), .Z(n333) );
  GTECH_XOR3 U355 ( .A(n346), .B(n358), .C(n356), .Z(n362) );
  GTECH_NAND2 U356 ( .A(I_a[5]), .B(I_b[0]), .Z(n356) );
  GTECH_OAI21 U357 ( .A(n363), .B(n364), .C(n365), .Z(n358) );
  GTECH_OAI21 U358 ( .A(n366), .B(n367), .C(n368), .Z(n365) );
  GTECH_NOT U359 ( .A(n369), .Z(n346) );
  GTECH_NAND2 U360 ( .A(I_a[4]), .B(I_b[1]), .Z(n369) );
  GTECH_ADD_ABC U361 ( .A(n370), .B(n371), .C(n372), .COUT(n341) );
  GTECH_XOR3 U362 ( .A(n366), .B(n368), .C(n363), .Z(n371) );
  GTECH_NOT U363 ( .A(n367), .Z(n363) );
  GTECH_OA21 U364 ( .A(n373), .B(n374), .C(n375), .Z(n370) );
  GTECH_XOR3 U365 ( .A(n351), .B(n353), .C(n352), .Z(n344) );
  GTECH_OAI21 U366 ( .A(n376), .B(n377), .C(n378), .Z(n352) );
  GTECH_NOT U367 ( .A(n379), .Z(n353) );
  GTECH_NAND2 U368 ( .A(I_b[3]), .B(I_a[2]), .Z(n379) );
  GTECH_NOT U369 ( .A(n349), .Z(n351) );
  GTECH_NAND2 U370 ( .A(I_b[2]), .B(I_a[3]), .Z(n349) );
  GTECH_NOT U371 ( .A(n380), .Z(n335) );
  GTECH_NAND3 U372 ( .A(I_a[0]), .B(n381), .C(I_b[4]), .Z(n380) );
  GTECH_NOT U373 ( .A(n382), .Z(n381) );
  GTECH_XNOR2 U374 ( .A(n383), .B(n382), .Z(N144) );
  GTECH_XOR3 U375 ( .A(n384), .B(n372), .C(n385), .Z(n382) );
  GTECH_OAI21 U376 ( .A(n373), .B(n374), .C(n375), .Z(n385) );
  GTECH_OAI21 U377 ( .A(n386), .B(n387), .C(n388), .Z(n375) );
  GTECH_NOT U378 ( .A(n373), .Z(n387) );
  GTECH_XOR3 U379 ( .A(n389), .B(n390), .C(n378), .Z(n372) );
  GTECH_NAND3 U380 ( .A(I_b[2]), .B(I_a[1]), .C(n391), .Z(n378) );
  GTECH_NOT U381 ( .A(n377), .Z(n390) );
  GTECH_NAND2 U382 ( .A(I_b[3]), .B(I_a[1]), .Z(n377) );
  GTECH_NOT U383 ( .A(n376), .Z(n389) );
  GTECH_NAND2 U384 ( .A(I_b[2]), .B(I_a[2]), .Z(n376) );
  GTECH_XOR3 U385 ( .A(n368), .B(n367), .C(n366), .Z(n384) );
  GTECH_NOT U386 ( .A(n364), .Z(n366) );
  GTECH_NAND2 U387 ( .A(I_a[4]), .B(I_b[0]), .Z(n364) );
  GTECH_OAI21 U388 ( .A(n392), .B(n393), .C(n394), .Z(n367) );
  GTECH_OAI21 U389 ( .A(n395), .B(n396), .C(n397), .Z(n394) );
  GTECH_NOT U390 ( .A(n396), .Z(n392) );
  GTECH_NOT U391 ( .A(n398), .Z(n368) );
  GTECH_NAND2 U392 ( .A(I_a[3]), .B(I_b[1]), .Z(n398) );
  GTECH_AND2 U393 ( .A(I_b[4]), .B(I_a[0]), .Z(n383) );
  GTECH_XOR3 U394 ( .A(n388), .B(n374), .C(n373), .Z(N143) );
  GTECH_XNOR2 U395 ( .A(n391), .B(n399), .Z(n373) );
  GTECH_AND2 U396 ( .A(I_b[2]), .B(I_a[1]), .Z(n399) );
  GTECH_NOT U397 ( .A(n400), .Z(n391) );
  GTECH_NAND2 U398 ( .A(I_b[3]), .B(I_a[0]), .Z(n400) );
  GTECH_NOT U399 ( .A(n386), .Z(n374) );
  GTECH_XOR3 U400 ( .A(n395), .B(n397), .C(n396), .Z(n386) );
  GTECH_OAI21 U401 ( .A(n401), .B(n402), .C(n403), .Z(n396) );
  GTECH_NOT U402 ( .A(n404), .Z(n397) );
  GTECH_NAND2 U403 ( .A(I_b[1]), .B(I_a[2]), .Z(n404) );
  GTECH_NOT U404 ( .A(n393), .Z(n395) );
  GTECH_NAND2 U405 ( .A(I_b[0]), .B(I_a[3]), .Z(n393) );
  GTECH_NOT U406 ( .A(n405), .Z(n388) );
  GTECH_NAND3 U407 ( .A(I_a[0]), .B(n406), .C(I_b[2]), .Z(n405) );
  GTECH_NOT U408 ( .A(n407), .Z(n406) );
  GTECH_XNOR2 U409 ( .A(n408), .B(n407), .Z(N142) );
  GTECH_XOR3 U410 ( .A(n409), .B(n410), .C(n403), .Z(n407) );
  GTECH_NAND3 U411 ( .A(n411), .B(I_b[0]), .C(I_a[1]), .Z(n403) );
  GTECH_NOT U412 ( .A(n401), .Z(n410) );
  GTECH_NAND2 U413 ( .A(I_a[1]), .B(I_b[1]), .Z(n401) );
  GTECH_NOT U414 ( .A(n402), .Z(n409) );
  GTECH_NAND2 U415 ( .A(I_b[0]), .B(I_a[2]), .Z(n402) );
  GTECH_AND2 U416 ( .A(I_b[2]), .B(I_a[0]), .Z(n408) );
  GTECH_XNOR2 U417 ( .A(n411), .B(n412), .Z(N141) );
  GTECH_NAND2 U418 ( .A(I_a[1]), .B(I_b[0]), .Z(n412) );
  GTECH_NOT U419 ( .A(n413), .Z(n411) );
  GTECH_NAND2 U420 ( .A(I_a[0]), .B(I_b[1]), .Z(n413) );
  GTECH_AND2 U421 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

