
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n113, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n113), .K(n113), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n250) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n113), .K(n113), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n113), .K(n113), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n113), .K(n113), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n113), .K(n113), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n113), .K(n113), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]) );
  GTECH_FJK1S A_reg_15_ ( .J(n113), .K(n113), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n266) );
  GTECH_FJK1S A_reg_14_ ( .J(n113), .K(n113), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n265) );
  GTECH_FJK1S A_reg_13_ ( .J(n113), .K(n113), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n264) );
  GTECH_FJK1S A_reg_12_ ( .J(n113), .K(n113), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n263) );
  GTECH_FJK1S A_reg_11_ ( .J(n113), .K(n113), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n262) );
  GTECH_FJK1S A_reg_10_ ( .J(n113), .K(n113), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n261) );
  GTECH_FJK1S A_reg_9_ ( .J(n113), .K(n113), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n260) );
  GTECH_FJK1S A_reg_8_ ( .J(n113), .K(n113), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n259) );
  GTECH_FJK1S A_reg_7_ ( .J(n113), .K(n113), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n258) );
  GTECH_FJK1S A_reg_6_ ( .J(n113), .K(n113), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n257) );
  GTECH_FJK1S A_reg_5_ ( .J(n113), .K(n113), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n256) );
  GTECH_FJK1S A_reg_4_ ( .J(n113), .K(n113), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n255) );
  GTECH_FJK1S A_reg_3_ ( .J(n113), .K(n113), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n254) );
  GTECH_FJK1S A_reg_2_ ( .J(n113), .K(n113), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n253) );
  GTECH_FJK1S A_reg_1_ ( .J(n113), .K(n113), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n252) );
  GTECH_FJK1S A_reg_0_ ( .J(n113), .K(n113), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n251) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n113), .K(n113), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n113), .K(n113), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n113), .K(n113), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n113), .K(n113), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n113), .K(n113), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n113), .K(n113), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n113), .K(n113), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n113), .K(n113), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n113), .K(n113), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n113), .K(n113), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n113), .K(n113), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n113), .K(n113), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n113), .K(n113), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n113), .K(n113), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n113), .K(n113), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n113), .K(n113), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n113), .K(n113), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n113), .K(n113), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n113), .K(n113), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n113), .K(n113), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n113), .K(n113), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n113), .K(n113), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n113), .K(n113), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n113), .K(n113), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n113), .K(n113), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n113), .K(n113), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n113), .K(n113), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n113), .K(n113), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n113), .K(n113), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n113), .K(n113), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n113), .K(n113), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n113), .K(n113), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n113), .K(n113), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n113), .K(n113), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n113), .K(n113), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n113), .K(n113), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n113), .K(n113), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n113), .K(n113), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n113), .K(n113), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n113), .K(n113), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n113), .K(n113), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n113), .K(n113), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n113), .K(n113), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n113), .K(n113), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n113), .K(n113), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n113), .K(n113), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n113), .K(n113), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n113), .K(n113), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n113), .K(n113), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n113), .K(n113), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n113), .K(n113), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n113), .K(n113), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n113), .K(n113), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n113), .K(n113), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n113), .K(n113), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n113), .K(n113), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n113), .K(n113), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n113), .K(n113), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n113), .K(n113), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n113), .K(n113), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n113), .K(n113), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n113), .K(n113), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n113), .K(n113), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n113), .K(n113), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n113), .K(n113), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n113), .K(n113), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U252 ( .Z(n113) );
  GTECH_NOT U253 ( .A(n268), .Z(N99) );
  GTECH_AOI222 U254 ( .A(n269), .B(n270), .C(n271), .D(n272), .E(n273), .F(
        n274), .Z(n268) );
  GTECH_NOT U255 ( .A(n275), .Z(N98) );
  GTECH_AOI222 U256 ( .A(n271), .B(n276), .C(n277), .D(n278), .E(R[15]), .F(
        n279), .Z(n275) );
  GTECH_NAND2 U257 ( .A(n280), .B(n281), .Z(n277) );
  GTECH_OAI2N2 U258 ( .A(n13), .B(n282), .C(R[14]), .D(n279), .Z(N97) );
  GTECH_OAI2N2 U259 ( .A(n14), .B(n282), .C(R[13]), .D(n279), .Z(N96) );
  GTECH_OAI2N2 U260 ( .A(n15), .B(n282), .C(R[12]), .D(n279), .Z(N95) );
  GTECH_OAI2N2 U261 ( .A(n16), .B(n282), .C(R[11]), .D(n279), .Z(N94) );
  GTECH_OAI2N2 U262 ( .A(n17), .B(n282), .C(R[10]), .D(n279), .Z(N93) );
  GTECH_OAI2N2 U263 ( .A(n18), .B(n282), .C(R[9]), .D(n279), .Z(N92) );
  GTECH_OAI2N2 U264 ( .A(n19), .B(n282), .C(R[8]), .D(n279), .Z(N91) );
  GTECH_OAI2N2 U265 ( .A(n20), .B(n282), .C(R[7]), .D(n279), .Z(N90) );
  GTECH_OAI2N2 U266 ( .A(n21), .B(n282), .C(R[6]), .D(n279), .Z(N89) );
  GTECH_OAI2N2 U267 ( .A(n22), .B(n282), .C(R[5]), .D(n279), .Z(N88) );
  GTECH_OAI2N2 U268 ( .A(n23), .B(n282), .C(R[4]), .D(n279), .Z(N87) );
  GTECH_OAI2N2 U269 ( .A(n24), .B(n282), .C(R[3]), .D(n279), .Z(N86) );
  GTECH_OAI2N2 U270 ( .A(n25), .B(n282), .C(R[2]), .D(n279), .Z(N85) );
  GTECH_OAI2N2 U271 ( .A(n26), .B(n282), .C(R[1]), .D(n279), .Z(N84) );
  GTECH_OAI2N2 U272 ( .A(n27), .B(n282), .C(R[0]), .D(n279), .Z(N83) );
  GTECH_AND2 U273 ( .A(M[15]), .B(n279), .Z(N42) );
  GTECH_AND2 U274 ( .A(M[14]), .B(n279), .Z(N39) );
  GTECH_AND2 U275 ( .A(M[13]), .B(n279), .Z(N38) );
  GTECH_AND2 U276 ( .A(M[12]), .B(n279), .Z(N37) );
  GTECH_AND2 U277 ( .A(M[11]), .B(n279), .Z(N36) );
  GTECH_AND2 U278 ( .A(M[10]), .B(n279), .Z(N35) );
  GTECH_AND2 U279 ( .A(M[9]), .B(n279), .Z(N34) );
  GTECH_AND2 U280 ( .A(M[8]), .B(n279), .Z(N33) );
  GTECH_AND2 U281 ( .A(M[7]), .B(n279), .Z(N32) );
  GTECH_AND2 U282 ( .A(M[6]), .B(n279), .Z(N31) );
  GTECH_AND2 U283 ( .A(M[5]), .B(n279), .Z(N30) );
  GTECH_AND2 U284 ( .A(M[4]), .B(n279), .Z(N29) );
  GTECH_AND2 U285 ( .A(M[3]), .B(n279), .Z(N28) );
  GTECH_AND2 U286 ( .A(M[2]), .B(n279), .Z(N27) );
  GTECH_AND2 U287 ( .A(M[1]), .B(n279), .Z(N26) );
  GTECH_AND2 U288 ( .A(M[0]), .B(n279), .Z(N25) );
  GTECH_NOT U289 ( .A(n283), .Z(n279) );
  GTECH_NAND2 U290 ( .A(n283), .B(n284), .Z(N19) );
  GTECH_NAND3 U291 ( .A(n285), .B(n286), .C(n287), .Z(n284) );
  GTECH_NAND3 U292 ( .A(n288), .B(n289), .C(n282), .Z(N18) );
  GTECH_AND2 U293 ( .A(n287), .B(n290), .Z(N17) );
  GTECH_OAI21 U294 ( .A(n8), .B(n291), .C(n285), .Z(n290) );
  GTECH_AND2 U295 ( .A(n287), .B(n292), .Z(N16) );
  GTECH_OAI21 U296 ( .A(n7), .B(n293), .C(n294), .Z(n292) );
  GTECH_NOT U297 ( .A(n295), .Z(N152) );
  GTECH_AOI222 U298 ( .A(n296), .B(n297), .C(n298), .D(n299), .E(n300), .F(
        n301), .Z(n295) );
  GTECH_NAND2 U299 ( .A(n289), .B(n302), .Z(N151) );
  GTECH_NOT U300 ( .A(n303), .Z(N150) );
  GTECH_AOI222 U301 ( .A(n304), .B(n296), .C(n298), .D(n305), .E(n300), .F(
        n306), .Z(n303) );
  GTECH_OAI21 U302 ( .A(n307), .B(n308), .C(n309), .Z(N15) );
  GTECH_NAND3 U303 ( .A(n287), .B(n310), .C(n307), .Z(n309) );
  GTECH_NOT U304 ( .A(n6), .Z(n307) );
  GTECH_NOT U305 ( .A(n311), .Z(N149) );
  GTECH_AOI222 U306 ( .A(n312), .B(n296), .C(n298), .D(n313), .E(n300), .F(
        n314), .Z(n311) );
  GTECH_NOT U307 ( .A(n315), .Z(N148) );
  GTECH_AOI222 U308 ( .A(n316), .B(n296), .C(n298), .D(n317), .E(n300), .F(
        n318), .Z(n315) );
  GTECH_NOT U309 ( .A(n319), .Z(N147) );
  GTECH_AOI222 U310 ( .A(n320), .B(n296), .C(n298), .D(n321), .E(n300), .F(
        n322), .Z(n319) );
  GTECH_NOT U311 ( .A(n323), .Z(N146) );
  GTECH_AOI222 U312 ( .A(n324), .B(n296), .C(n298), .D(n325), .E(n300), .F(
        n326), .Z(n323) );
  GTECH_NOT U313 ( .A(n327), .Z(N145) );
  GTECH_AOI222 U314 ( .A(n328), .B(n296), .C(n298), .D(n329), .E(n300), .F(
        n330), .Z(n327) );
  GTECH_NOT U315 ( .A(n331), .Z(N144) );
  GTECH_AOI222 U316 ( .A(n332), .B(n296), .C(n298), .D(n333), .E(n300), .F(
        n334), .Z(n331) );
  GTECH_NOT U317 ( .A(n335), .Z(N143) );
  GTECH_AOI222 U318 ( .A(n336), .B(n296), .C(n298), .D(n337), .E(n300), .F(
        n338), .Z(n335) );
  GTECH_NOT U319 ( .A(n339), .Z(N142) );
  GTECH_AOI222 U320 ( .A(n340), .B(n296), .C(n298), .D(n341), .E(n300), .F(
        n342), .Z(n339) );
  GTECH_NOT U321 ( .A(n343), .Z(N141) );
  GTECH_AOI222 U322 ( .A(n344), .B(n296), .C(n298), .D(n345), .E(n300), .F(
        n346), .Z(n343) );
  GTECH_NOT U323 ( .A(n347), .Z(N140) );
  GTECH_AOI222 U324 ( .A(n348), .B(n296), .C(n298), .D(n349), .E(n300), .F(
        n350), .Z(n347) );
  GTECH_NOT U325 ( .A(n308), .Z(N14) );
  GTECH_NAND2 U326 ( .A(n287), .B(n250), .Z(n308) );
  GTECH_NOT U327 ( .A(n351), .Z(N139) );
  GTECH_AOI222 U328 ( .A(n352), .B(n296), .C(n298), .D(n353), .E(n300), .F(
        n354), .Z(n351) );
  GTECH_NOT U329 ( .A(n355), .Z(N138) );
  GTECH_AOI222 U330 ( .A(n356), .B(n296), .C(n298), .D(n357), .E(n300), .F(
        n358), .Z(n355) );
  GTECH_NOT U331 ( .A(n359), .Z(N137) );
  GTECH_AOI222 U332 ( .A(n360), .B(n296), .C(n298), .D(n361), .E(n300), .F(
        n362), .Z(n359) );
  GTECH_NOT U333 ( .A(n363), .Z(N136) );
  GTECH_AOI222 U334 ( .A(n296), .B(n270), .C(n298), .D(n272), .E(n300), .F(
        n274), .Z(n363) );
  GTECH_NOT U335 ( .A(n364), .Z(n274) );
  GTECH_XOR2 U336 ( .A(n365), .B(n366), .Z(n364) );
  GTECH_NOT U337 ( .A(n367), .Z(n366) );
  GTECH_NOT U338 ( .A(n368), .Z(n298) );
  GTECH_NOT U339 ( .A(n369), .Z(n270) );
  GTECH_XOR2 U340 ( .A(n365), .B(n370), .Z(n369) );
  GTECH_NOT U341 ( .A(n371), .Z(n370) );
  GTECH_XOR2 U342 ( .A(n272), .B(n252), .Z(n365) );
  GTECH_OAI21 U343 ( .A(n12), .B(n368), .C(n372), .Z(N135) );
  GTECH_OAI21 U344 ( .A(n300), .B(n296), .C(n278), .Z(n372) );
  GTECH_OAI21 U345 ( .A(n12), .B(n373), .C(n367), .Z(n278) );
  GTECH_NOT U346 ( .A(n374), .Z(n296) );
  GTECH_NAND3 U347 ( .A(n28), .B(n375), .C(N155), .Z(n374) );
  GTECH_NOT U348 ( .A(n376), .Z(n300) );
  GTECH_NAND3 U349 ( .A(n10), .B(n377), .C(N155), .Z(n376) );
  GTECH_NAND2 U350 ( .A(n378), .B(N155), .Z(n368) );
  GTECH_XOR2 U351 ( .A(n375), .B(n28), .Z(n378) );
  GTECH_AND2 U352 ( .A(N155), .B(n379), .Z(N134) );
  GTECH_NOT U353 ( .A(n13), .Z(n379) );
  GTECH_AND2 U354 ( .A(N155), .B(n380), .Z(N133) );
  GTECH_NOT U355 ( .A(n14), .Z(n380) );
  GTECH_AND2 U356 ( .A(N155), .B(n381), .Z(N132) );
  GTECH_NOT U357 ( .A(n15), .Z(n381) );
  GTECH_AND2 U358 ( .A(N155), .B(n382), .Z(N131) );
  GTECH_NOT U359 ( .A(n16), .Z(n382) );
  GTECH_AND2 U360 ( .A(N155), .B(n383), .Z(N130) );
  GTECH_NOT U361 ( .A(n17), .Z(n383) );
  GTECH_AND2 U362 ( .A(N155), .B(n384), .Z(N129) );
  GTECH_NOT U363 ( .A(n18), .Z(n384) );
  GTECH_AND2 U364 ( .A(N155), .B(n385), .Z(N128) );
  GTECH_NOT U365 ( .A(n19), .Z(n385) );
  GTECH_AND2 U366 ( .A(N155), .B(n386), .Z(N127) );
  GTECH_NOT U367 ( .A(n20), .Z(n386) );
  GTECH_AND2 U368 ( .A(N155), .B(n387), .Z(N126) );
  GTECH_NOT U369 ( .A(n21), .Z(n387) );
  GTECH_AND2 U370 ( .A(N155), .B(n388), .Z(N125) );
  GTECH_NOT U371 ( .A(n22), .Z(n388) );
  GTECH_AND2 U372 ( .A(N155), .B(n389), .Z(N124) );
  GTECH_NOT U373 ( .A(n23), .Z(n389) );
  GTECH_AND2 U374 ( .A(N155), .B(n390), .Z(N123) );
  GTECH_NOT U375 ( .A(n24), .Z(n390) );
  GTECH_AND2 U376 ( .A(N155), .B(n391), .Z(N122) );
  GTECH_NOT U377 ( .A(n25), .Z(n391) );
  GTECH_AND2 U378 ( .A(N155), .B(n392), .Z(N121) );
  GTECH_NOT U379 ( .A(n26), .Z(n392) );
  GTECH_AND2 U380 ( .A(N155), .B(n393), .Z(N120) );
  GTECH_NOT U381 ( .A(n27), .Z(n393) );
  GTECH_NOT U382 ( .A(n302), .Z(N155) );
  GTECH_NAND3 U383 ( .A(n7), .B(n8), .C(n394), .Z(n302) );
  GTECH_AND4 U384 ( .A(n310), .B(n6), .C(n289), .D(n9), .Z(n394) );
  GTECH_NOT U385 ( .A(n250), .Z(n310) );
  GTECH_NOT U386 ( .A(n395), .Z(N116) );
  GTECH_AOI222 U387 ( .A(n271), .B(n299), .C(n273), .D(n301), .E(n297), .F(
        n269), .Z(n395) );
  GTECH_XOR2 U388 ( .A(n396), .B(n397), .Z(n297) );
  GTECH_ADD_ABC U389 ( .A(n31), .B(n266), .C(n398), .COUT(n397) );
  GTECH_XOR2 U390 ( .A(n399), .B(n396), .Z(n301) );
  GTECH_XOR2 U391 ( .A(A[16]), .B(n30), .Z(n396) );
  GTECH_OAI21 U392 ( .A(n400), .B(n31), .C(n401), .Z(n399) );
  GTECH_OAI21 U393 ( .A(n266), .B(n305), .C(n402), .Z(n401) );
  GTECH_NOT U394 ( .A(n30), .Z(n299) );
  GTECH_NAND2 U395 ( .A(n282), .B(n403), .Z(N115) );
  GTECH_NOT U396 ( .A(N41), .Z(n403) );
  GTECH_NAND2 U397 ( .A(n289), .B(n283), .Z(N41) );
  GTECH_NAND2 U398 ( .A(Ld), .B(n289), .Z(n283) );
  GTECH_NOT U399 ( .A(n404), .Z(N113) );
  GTECH_AOI222 U400 ( .A(n271), .B(n305), .C(n273), .D(n306), .E(n304), .F(
        n269), .Z(n404) );
  GTECH_XOR2 U401 ( .A(n405), .B(n398), .Z(n304) );
  GTECH_ADD_ABC U402 ( .A(n32), .B(n265), .C(n406), .COUT(n398) );
  GTECH_NOT U403 ( .A(n407), .Z(n306) );
  GTECH_XOR2 U404 ( .A(n405), .B(n408), .Z(n407) );
  GTECH_NOT U405 ( .A(n402), .Z(n408) );
  GTECH_OAI21 U406 ( .A(n32), .B(n409), .C(n410), .Z(n402) );
  GTECH_OAI21 U407 ( .A(n265), .B(n313), .C(n411), .Z(n410) );
  GTECH_XOR2 U408 ( .A(n400), .B(n31), .Z(n405) );
  GTECH_NOT U409 ( .A(n266), .Z(n400) );
  GTECH_NOT U410 ( .A(n31), .Z(n305) );
  GTECH_NOT U411 ( .A(n412), .Z(N112) );
  GTECH_AOI222 U412 ( .A(n271), .B(n313), .C(n273), .D(n314), .E(n312), .F(
        n269), .Z(n412) );
  GTECH_XOR2 U413 ( .A(n413), .B(n406), .Z(n312) );
  GTECH_ADD_ABC U414 ( .A(n33), .B(n264), .C(n414), .COUT(n406) );
  GTECH_NOT U415 ( .A(n415), .Z(n314) );
  GTECH_XOR2 U416 ( .A(n413), .B(n416), .Z(n415) );
  GTECH_NOT U417 ( .A(n411), .Z(n416) );
  GTECH_OAI21 U418 ( .A(n33), .B(n417), .C(n418), .Z(n411) );
  GTECH_OAI21 U419 ( .A(n264), .B(n317), .C(n419), .Z(n418) );
  GTECH_XOR2 U420 ( .A(n409), .B(n32), .Z(n413) );
  GTECH_NOT U421 ( .A(n265), .Z(n409) );
  GTECH_NOT U422 ( .A(n32), .Z(n313) );
  GTECH_NOT U423 ( .A(n420), .Z(N111) );
  GTECH_AOI222 U424 ( .A(n271), .B(n317), .C(n273), .D(n318), .E(n316), .F(
        n269), .Z(n420) );
  GTECH_XOR2 U425 ( .A(n421), .B(n414), .Z(n316) );
  GTECH_ADD_ABC U426 ( .A(n34), .B(n263), .C(n422), .COUT(n414) );
  GTECH_NOT U427 ( .A(n423), .Z(n318) );
  GTECH_XOR2 U428 ( .A(n421), .B(n424), .Z(n423) );
  GTECH_NOT U429 ( .A(n419), .Z(n424) );
  GTECH_OAI21 U430 ( .A(n34), .B(n425), .C(n426), .Z(n419) );
  GTECH_OAI21 U431 ( .A(n263), .B(n321), .C(n427), .Z(n426) );
  GTECH_XOR2 U432 ( .A(n417), .B(n33), .Z(n421) );
  GTECH_NOT U433 ( .A(n264), .Z(n417) );
  GTECH_NOT U434 ( .A(n33), .Z(n317) );
  GTECH_NOT U435 ( .A(n428), .Z(N110) );
  GTECH_AOI222 U436 ( .A(n271), .B(n321), .C(n273), .D(n322), .E(n320), .F(
        n269), .Z(n428) );
  GTECH_XOR2 U437 ( .A(n429), .B(n422), .Z(n320) );
  GTECH_ADD_ABC U438 ( .A(n35), .B(n262), .C(n430), .COUT(n422) );
  GTECH_NOT U439 ( .A(n431), .Z(n322) );
  GTECH_XOR2 U440 ( .A(n429), .B(n432), .Z(n431) );
  GTECH_NOT U441 ( .A(n427), .Z(n432) );
  GTECH_OAI21 U442 ( .A(n35), .B(n433), .C(n434), .Z(n427) );
  GTECH_OAI21 U443 ( .A(n262), .B(n325), .C(n435), .Z(n434) );
  GTECH_XOR2 U444 ( .A(n425), .B(n34), .Z(n429) );
  GTECH_NOT U445 ( .A(n263), .Z(n425) );
  GTECH_NOT U446 ( .A(n34), .Z(n321) );
  GTECH_NOT U447 ( .A(n436), .Z(N109) );
  GTECH_AOI222 U448 ( .A(n271), .B(n325), .C(n273), .D(n326), .E(n324), .F(
        n269), .Z(n436) );
  GTECH_XOR2 U449 ( .A(n437), .B(n430), .Z(n324) );
  GTECH_ADD_ABC U450 ( .A(n36), .B(n261), .C(n438), .COUT(n430) );
  GTECH_NOT U451 ( .A(n439), .Z(n326) );
  GTECH_XOR2 U452 ( .A(n437), .B(n440), .Z(n439) );
  GTECH_NOT U453 ( .A(n435), .Z(n440) );
  GTECH_OAI21 U454 ( .A(n36), .B(n441), .C(n442), .Z(n435) );
  GTECH_OAI21 U455 ( .A(n261), .B(n329), .C(n443), .Z(n442) );
  GTECH_XOR2 U456 ( .A(n433), .B(n35), .Z(n437) );
  GTECH_NOT U457 ( .A(n262), .Z(n433) );
  GTECH_NOT U458 ( .A(n35), .Z(n325) );
  GTECH_NOT U459 ( .A(n444), .Z(N108) );
  GTECH_AOI222 U460 ( .A(n271), .B(n329), .C(n273), .D(n330), .E(n328), .F(
        n269), .Z(n444) );
  GTECH_XOR2 U461 ( .A(n445), .B(n438), .Z(n328) );
  GTECH_ADD_ABC U462 ( .A(n37), .B(n260), .C(n446), .COUT(n438) );
  GTECH_NOT U463 ( .A(n447), .Z(n330) );
  GTECH_XOR2 U464 ( .A(n445), .B(n448), .Z(n447) );
  GTECH_NOT U465 ( .A(n443), .Z(n448) );
  GTECH_OAI21 U466 ( .A(n37), .B(n449), .C(n450), .Z(n443) );
  GTECH_OAI21 U467 ( .A(n260), .B(n333), .C(n451), .Z(n450) );
  GTECH_XOR2 U468 ( .A(n441), .B(n36), .Z(n445) );
  GTECH_NOT U469 ( .A(n261), .Z(n441) );
  GTECH_NOT U470 ( .A(n36), .Z(n329) );
  GTECH_NOT U471 ( .A(n452), .Z(N107) );
  GTECH_AOI222 U472 ( .A(n271), .B(n333), .C(n273), .D(n334), .E(n332), .F(
        n269), .Z(n452) );
  GTECH_XOR2 U473 ( .A(n453), .B(n446), .Z(n332) );
  GTECH_ADD_ABC U474 ( .A(n38), .B(n259), .C(n454), .COUT(n446) );
  GTECH_NOT U475 ( .A(n455), .Z(n334) );
  GTECH_XOR2 U476 ( .A(n453), .B(n456), .Z(n455) );
  GTECH_NOT U477 ( .A(n451), .Z(n456) );
  GTECH_OAI21 U478 ( .A(n38), .B(n457), .C(n458), .Z(n451) );
  GTECH_OAI21 U479 ( .A(n259), .B(n337), .C(n459), .Z(n458) );
  GTECH_XOR2 U480 ( .A(n449), .B(n37), .Z(n453) );
  GTECH_NOT U481 ( .A(n260), .Z(n449) );
  GTECH_NOT U482 ( .A(n37), .Z(n333) );
  GTECH_NOT U483 ( .A(n460), .Z(N106) );
  GTECH_AOI222 U484 ( .A(n271), .B(n337), .C(n273), .D(n338), .E(n336), .F(
        n269), .Z(n460) );
  GTECH_XOR2 U485 ( .A(n461), .B(n454), .Z(n336) );
  GTECH_ADD_ABC U486 ( .A(n39), .B(n258), .C(n462), .COUT(n454) );
  GTECH_NOT U487 ( .A(n463), .Z(n338) );
  GTECH_XOR2 U488 ( .A(n461), .B(n464), .Z(n463) );
  GTECH_NOT U489 ( .A(n459), .Z(n464) );
  GTECH_OAI21 U490 ( .A(n39), .B(n465), .C(n466), .Z(n459) );
  GTECH_OAI21 U491 ( .A(n258), .B(n341), .C(n467), .Z(n466) );
  GTECH_XOR2 U492 ( .A(n457), .B(n38), .Z(n461) );
  GTECH_NOT U493 ( .A(n259), .Z(n457) );
  GTECH_NOT U494 ( .A(n38), .Z(n337) );
  GTECH_NOT U495 ( .A(n468), .Z(N105) );
  GTECH_AOI222 U496 ( .A(n271), .B(n341), .C(n273), .D(n342), .E(n340), .F(
        n269), .Z(n468) );
  GTECH_XOR2 U497 ( .A(n469), .B(n462), .Z(n340) );
  GTECH_ADD_ABC U498 ( .A(n40), .B(n257), .C(n470), .COUT(n462) );
  GTECH_NOT U499 ( .A(n471), .Z(n342) );
  GTECH_XOR2 U500 ( .A(n469), .B(n472), .Z(n471) );
  GTECH_NOT U501 ( .A(n467), .Z(n472) );
  GTECH_OAI21 U502 ( .A(n40), .B(n473), .C(n474), .Z(n467) );
  GTECH_OAI21 U503 ( .A(n257), .B(n345), .C(n475), .Z(n474) );
  GTECH_XOR2 U504 ( .A(n465), .B(n39), .Z(n469) );
  GTECH_NOT U505 ( .A(n258), .Z(n465) );
  GTECH_NOT U506 ( .A(n39), .Z(n341) );
  GTECH_NOT U507 ( .A(n476), .Z(N104) );
  GTECH_AOI222 U508 ( .A(n271), .B(n345), .C(n273), .D(n346), .E(n344), .F(
        n269), .Z(n476) );
  GTECH_XOR2 U509 ( .A(n477), .B(n470), .Z(n344) );
  GTECH_ADD_ABC U510 ( .A(n41), .B(n256), .C(n478), .COUT(n470) );
  GTECH_NOT U511 ( .A(n479), .Z(n346) );
  GTECH_XOR2 U512 ( .A(n477), .B(n480), .Z(n479) );
  GTECH_NOT U513 ( .A(n475), .Z(n480) );
  GTECH_OAI21 U514 ( .A(n41), .B(n481), .C(n482), .Z(n475) );
  GTECH_OAI21 U515 ( .A(n256), .B(n349), .C(n483), .Z(n482) );
  GTECH_XOR2 U516 ( .A(n473), .B(n40), .Z(n477) );
  GTECH_NOT U517 ( .A(n257), .Z(n473) );
  GTECH_NOT U518 ( .A(n40), .Z(n345) );
  GTECH_NOT U519 ( .A(n484), .Z(N103) );
  GTECH_AOI222 U520 ( .A(n271), .B(n349), .C(n273), .D(n350), .E(n348), .F(
        n269), .Z(n484) );
  GTECH_XOR2 U521 ( .A(n485), .B(n478), .Z(n348) );
  GTECH_ADD_ABC U522 ( .A(n42), .B(n255), .C(n486), .COUT(n478) );
  GTECH_NOT U523 ( .A(n487), .Z(n350) );
  GTECH_XOR2 U524 ( .A(n485), .B(n488), .Z(n487) );
  GTECH_NOT U525 ( .A(n483), .Z(n488) );
  GTECH_OAI21 U526 ( .A(n42), .B(n489), .C(n490), .Z(n483) );
  GTECH_OAI21 U527 ( .A(n255), .B(n353), .C(n491), .Z(n490) );
  GTECH_XOR2 U528 ( .A(n481), .B(n41), .Z(n485) );
  GTECH_NOT U529 ( .A(n256), .Z(n481) );
  GTECH_NOT U530 ( .A(n41), .Z(n349) );
  GTECH_NOT U531 ( .A(n492), .Z(N102) );
  GTECH_AOI222 U532 ( .A(n271), .B(n353), .C(n273), .D(n354), .E(n352), .F(
        n269), .Z(n492) );
  GTECH_XOR2 U533 ( .A(n493), .B(n486), .Z(n352) );
  GTECH_ADD_ABC U534 ( .A(n43), .B(n254), .C(n494), .COUT(n486) );
  GTECH_NOT U535 ( .A(n495), .Z(n354) );
  GTECH_XOR2 U536 ( .A(n493), .B(n496), .Z(n495) );
  GTECH_NOT U537 ( .A(n491), .Z(n496) );
  GTECH_OAI21 U538 ( .A(n43), .B(n497), .C(n498), .Z(n491) );
  GTECH_OAI21 U539 ( .A(n254), .B(n357), .C(n499), .Z(n498) );
  GTECH_XOR2 U540 ( .A(n489), .B(n42), .Z(n493) );
  GTECH_NOT U541 ( .A(n255), .Z(n489) );
  GTECH_NOT U542 ( .A(n42), .Z(n353) );
  GTECH_NOT U543 ( .A(n500), .Z(N101) );
  GTECH_AOI222 U544 ( .A(n271), .B(n357), .C(n273), .D(n358), .E(n356), .F(
        n269), .Z(n500) );
  GTECH_XOR2 U545 ( .A(n501), .B(n494), .Z(n356) );
  GTECH_ADD_ABC U546 ( .A(n29), .B(n253), .C(n502), .COUT(n494) );
  GTECH_NOT U547 ( .A(n503), .Z(n358) );
  GTECH_XOR2 U548 ( .A(n501), .B(n504), .Z(n503) );
  GTECH_NOT U549 ( .A(n499), .Z(n504) );
  GTECH_OAI21 U550 ( .A(n29), .B(n505), .C(n506), .Z(n499) );
  GTECH_OAI21 U551 ( .A(n253), .B(n361), .C(n507), .Z(n506) );
  GTECH_XOR2 U552 ( .A(n497), .B(n43), .Z(n501) );
  GTECH_NOT U553 ( .A(n254), .Z(n497) );
  GTECH_NOT U554 ( .A(n43), .Z(n357) );
  GTECH_NOT U555 ( .A(n508), .Z(N100) );
  GTECH_AOI222 U556 ( .A(n360), .B(n269), .C(n271), .D(n361), .E(n273), .F(
        n362), .Z(n508) );
  GTECH_NOT U557 ( .A(n509), .Z(n362) );
  GTECH_XOR2 U558 ( .A(n510), .B(n511), .Z(n509) );
  GTECH_NOT U559 ( .A(n507), .Z(n511) );
  GTECH_OAI21 U560 ( .A(n11), .B(n512), .C(n513), .Z(n507) );
  GTECH_OAI21 U561 ( .A(n252), .B(n272), .C(n367), .Z(n513) );
  GTECH_NAND2 U562 ( .A(n12), .B(n373), .Z(n367) );
  GTECH_NOT U563 ( .A(n11), .Z(n272) );
  GTECH_NOT U564 ( .A(n252), .Z(n512) );
  GTECH_NOT U565 ( .A(n281), .Z(n273) );
  GTECH_NAND2 U566 ( .A(N82), .B(n10), .Z(n281) );
  GTECH_NOT U567 ( .A(n514), .Z(N82) );
  GTECH_NOT U568 ( .A(n29), .Z(n361) );
  GTECH_OAI21 U569 ( .A(n10), .B(n514), .C(n515), .Z(n271) );
  GTECH_NAND3 U570 ( .A(n28), .B(n287), .C(n10), .Z(n515) );
  GTECH_NAND2 U571 ( .A(n287), .B(n377), .Z(n514) );
  GTECH_NOT U572 ( .A(n28), .Z(n377) );
  GTECH_NOT U573 ( .A(n280), .Z(n269) );
  GTECH_NAND3 U574 ( .A(n287), .B(n375), .C(n28), .Z(n280) );
  GTECH_NOT U575 ( .A(n10), .Z(n375) );
  GTECH_NOT U576 ( .A(n282), .Z(n287) );
  GTECH_OAI21 U577 ( .A(n285), .B(n286), .C(n516), .Z(n282) );
  GTECH_AND2 U578 ( .A(n288), .B(n289), .Z(n516) );
  GTECH_NOT U579 ( .A(Rst), .Z(n289) );
  GTECH_NOT U580 ( .A(Ld), .Z(n288) );
  GTECH_NOT U581 ( .A(n9), .Z(n286) );
  GTECH_NAND2 U582 ( .A(n8), .B(n291), .Z(n285) );
  GTECH_NOT U583 ( .A(n294), .Z(n291) );
  GTECH_NAND2 U584 ( .A(n7), .B(n293), .Z(n294) );
  GTECH_NOT U585 ( .A(n517), .Z(n293) );
  GTECH_NAND2 U586 ( .A(n6), .B(n250), .Z(n517) );
  GTECH_XOR2 U587 ( .A(n510), .B(n502), .Z(n360) );
  GTECH_ADD_ABC U588 ( .A(n252), .B(n11), .C(n371), .COUT(n502) );
  GTECH_NAND2 U589 ( .A(n276), .B(n373), .Z(n371) );
  GTECH_NOT U590 ( .A(n251), .Z(n373) );
  GTECH_NOT U591 ( .A(n12), .Z(n276) );
  GTECH_XOR2 U592 ( .A(n505), .B(n29), .Z(n510) );
  GTECH_NOT U593 ( .A(n253), .Z(n505) );
endmodule

