
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378;

  GTECH_MUX2 U131 ( .A(n270), .B(n271), .S(n272), .Z(sum[9]) );
  GTECH_XNOR2 U132 ( .A(n273), .B(n274), .Z(n271) );
  GTECH_XOR2 U133 ( .A(n275), .B(n274), .Z(n270) );
  GTECH_OAI21 U134 ( .A(a[9]), .B(b[9]), .C(n276), .Z(n274) );
  GTECH_NAND2 U135 ( .A(n277), .B(n278), .Z(sum[8]) );
  GTECH_OAI21 U136 ( .A(n273), .B(n275), .C(n279), .Z(n277) );
  GTECH_MUX2 U137 ( .A(n280), .B(n281), .S(n282), .Z(sum[7]) );
  GTECH_XNOR2 U138 ( .A(n283), .B(n284), .Z(n281) );
  GTECH_XOR2 U139 ( .A(n283), .B(n285), .Z(n280) );
  GTECH_OA21 U140 ( .A(n286), .B(n287), .C(n288), .Z(n285) );
  GTECH_NOR2 U141 ( .A(b[6]), .B(a[6]), .Z(n286) );
  GTECH_XNOR2 U142 ( .A(a[7]), .B(b[7]), .Z(n283) );
  GTECH_MUX2 U143 ( .A(n289), .B(n290), .S(n282), .Z(sum[6]) );
  GTECH_XNOR2 U144 ( .A(n291), .B(n292), .Z(n290) );
  GTECH_XOR2 U145 ( .A(n291), .B(n287), .Z(n289) );
  GTECH_ADD_AB U146 ( .A(n293), .B(n294), .COUT(n287) );
  GTECH_OAI21 U147 ( .A(b[5]), .B(a[5]), .C(n295), .Z(n293) );
  GTECH_OAI21 U148 ( .A(b[6]), .B(a[6]), .C(n288), .Z(n291) );
  GTECH_MUX2 U149 ( .A(n296), .B(n297), .S(n298), .Z(sum[5]) );
  GTECH_OA21 U150 ( .A(b[5]), .B(a[5]), .C(n294), .Z(n298) );
  GTECH_OAI21 U151 ( .A(n295), .B(n282), .C(n299), .Z(n297) );
  GTECH_NOT U152 ( .A(n300), .Z(n296) );
  GTECH_AOI21 U153 ( .A(n299), .B(n282), .C(n295), .Z(n300) );
  GTECH_AND_NOT U154 ( .A(a[4]), .B(n301), .Z(n295) );
  GTECH_XNOR2 U155 ( .A(n302), .B(n282), .Z(sum[4]) );
  GTECH_MUX2 U156 ( .A(n303), .B(n304), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U157 ( .A(n305), .B(n306), .Z(n304) );
  GTECH_XNOR2 U158 ( .A(n305), .B(n307), .Z(n303) );
  GTECH_OA21 U159 ( .A(n308), .B(n309), .C(n310), .Z(n307) );
  GTECH_XOR2 U160 ( .A(a[3]), .B(b[3]), .Z(n305) );
  GTECH_MUX2 U161 ( .A(n311), .B(n312), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U162 ( .A(n313), .B(n314), .Z(n312) );
  GTECH_XOR2 U163 ( .A(n309), .B(n313), .Z(n311) );
  GTECH_OR_NOT U164 ( .A(n308), .B(n310), .Z(n313) );
  GTECH_OA21 U165 ( .A(n315), .B(n316), .C(n317), .Z(n309) );
  GTECH_MUX2 U166 ( .A(n318), .B(n319), .S(n320), .Z(sum[1]) );
  GTECH_AND_NOT U167 ( .A(n317), .B(n315), .Z(n320) );
  GTECH_NOT U168 ( .A(n321), .Z(n319) );
  GTECH_AOI21 U169 ( .A(n322), .B(n316), .C(n323), .Z(n321) );
  GTECH_OAI21 U170 ( .A(n323), .B(n322), .C(n316), .Z(n318) );
  GTECH_MUX2 U171 ( .A(n324), .B(n325), .S(n326), .Z(sum[15]) );
  GTECH_XOR2 U172 ( .A(n327), .B(n328), .Z(n325) );
  GTECH_XNOR2 U173 ( .A(n327), .B(n329), .Z(n324) );
  GTECH_AOI21 U174 ( .A(n330), .B(n331), .C(n332), .Z(n329) );
  GTECH_OR2 U175 ( .A(b[14]), .B(a[14]), .Z(n330) );
  GTECH_XOR2 U176 ( .A(a[15]), .B(b[15]), .Z(n327) );
  GTECH_MUX2 U177 ( .A(n333), .B(n334), .S(n326), .Z(sum[14]) );
  GTECH_XNOR2 U178 ( .A(n335), .B(n336), .Z(n334) );
  GTECH_XNOR2 U179 ( .A(n331), .B(n336), .Z(n333) );
  GTECH_OAI21 U180 ( .A(b[14]), .B(a[14]), .C(n337), .Z(n336) );
  GTECH_AOI21 U181 ( .A(n338), .B(n339), .C(n340), .Z(n331) );
  GTECH_MUX2 U182 ( .A(n341), .B(n342), .S(n326), .Z(sum[13]) );
  GTECH_XNOR2 U183 ( .A(n343), .B(n344), .Z(n342) );
  GTECH_XOR2 U184 ( .A(n345), .B(n343), .Z(n341) );
  GTECH_OA21 U185 ( .A(a[13]), .B(b[13]), .C(n338), .Z(n343) );
  GTECH_NAND2 U186 ( .A(n346), .B(n347), .Z(sum[12]) );
  GTECH_OAI21 U187 ( .A(n345), .B(n344), .C(n326), .Z(n346) );
  GTECH_MUX2 U188 ( .A(n348), .B(n349), .S(n272), .Z(sum[11]) );
  GTECH_XOR2 U189 ( .A(n350), .B(n351), .Z(n349) );
  GTECH_OA21 U190 ( .A(n352), .B(n353), .C(n354), .Z(n351) );
  GTECH_NOT U191 ( .A(n355), .Z(n353) );
  GTECH_XNOR2 U192 ( .A(n350), .B(n356), .Z(n348) );
  GTECH_XNOR2 U193 ( .A(a[11]), .B(b[11]), .Z(n350) );
  GTECH_MUX2 U194 ( .A(n357), .B(n358), .S(n272), .Z(sum[10]) );
  GTECH_XNOR2 U195 ( .A(n359), .B(n355), .Z(n358) );
  GTECH_AOI21 U196 ( .A(n276), .B(n360), .C(n361), .Z(n355) );
  GTECH_XOR2 U197 ( .A(n359), .B(n362), .Z(n357) );
  GTECH_OR_NOT U198 ( .A(n352), .B(n354), .Z(n359) );
  GTECH_XNOR2 U199 ( .A(n322), .B(n363), .Z(sum[0]) );
  GTECH_NOT U200 ( .A(cin), .Z(n322) );
  GTECH_OAI21 U201 ( .A(n364), .B(n365), .C(n347), .Z(cout) );
  GTECH_OR3 U202 ( .A(n345), .B(n344), .C(n326), .Z(n347) );
  GTECH_NOT U203 ( .A(n364), .Z(n326) );
  GTECH_NOT U204 ( .A(n339), .Z(n345) );
  GTECH_NAND2 U205 ( .A(a[12]), .B(b[12]), .Z(n339) );
  GTECH_AOI21 U206 ( .A(n328), .B(a[15]), .C(n366), .Z(n365) );
  GTECH_OA21 U207 ( .A(a[15]), .B(n328), .C(b[15]), .Z(n366) );
  GTECH_NAND2 U208 ( .A(n337), .B(n367), .Z(n328) );
  GTECH_OAI21 U209 ( .A(a[14]), .B(b[14]), .C(n335), .Z(n367) );
  GTECH_AOI21 U210 ( .A(n338), .B(n344), .C(n340), .Z(n335) );
  GTECH_NOR2 U211 ( .A(b[13]), .B(a[13]), .Z(n340) );
  GTECH_NOR2 U212 ( .A(b[12]), .B(a[12]), .Z(n344) );
  GTECH_NAND2 U213 ( .A(a[13]), .B(b[13]), .Z(n338) );
  GTECH_NOT U214 ( .A(n332), .Z(n337) );
  GTECH_ADD_AB U215 ( .A(b[14]), .B(a[14]), .COUT(n332) );
  GTECH_OA21 U216 ( .A(n368), .B(n272), .C(n278), .Z(n364) );
  GTECH_OR3 U217 ( .A(n275), .B(n273), .C(n279), .Z(n278) );
  GTECH_NOT U218 ( .A(n272), .Z(n279) );
  GTECH_NOT U219 ( .A(n360), .Z(n273) );
  GTECH_NAND2 U220 ( .A(b[8]), .B(a[8]), .Z(n360) );
  GTECH_MUX2 U221 ( .A(n302), .B(n369), .S(n282), .Z(n272) );
  GTECH_MUX2 U222 ( .A(n363), .B(n370), .S(cin), .Z(n282) );
  GTECH_OA21 U223 ( .A(a[3]), .B(n306), .C(n371), .Z(n370) );
  GTECH_NOT U224 ( .A(n372), .Z(n371) );
  GTECH_AOI21 U225 ( .A(n306), .B(a[3]), .C(b[3]), .Z(n372) );
  GTECH_OAI21 U226 ( .A(n314), .B(n308), .C(n310), .Z(n306) );
  GTECH_NAND2 U227 ( .A(b[2]), .B(a[2]), .Z(n310) );
  GTECH_NOR2 U228 ( .A(a[2]), .B(b[2]), .Z(n308) );
  GTECH_OA21 U229 ( .A(n323), .B(n315), .C(n317), .Z(n314) );
  GTECH_NAND2 U230 ( .A(a[1]), .B(b[1]), .Z(n317) );
  GTECH_NOR2 U231 ( .A(b[1]), .B(a[1]), .Z(n315) );
  GTECH_AND_NOT U232 ( .A(n316), .B(n323), .Z(n363) );
  GTECH_NOR2 U233 ( .A(b[0]), .B(a[0]), .Z(n323) );
  GTECH_NAND2 U234 ( .A(a[0]), .B(b[0]), .Z(n316) );
  GTECH_AOI21 U235 ( .A(n284), .B(a[7]), .C(n373), .Z(n369) );
  GTECH_OA21 U236 ( .A(a[7]), .B(n284), .C(b[7]), .Z(n373) );
  GTECH_NAND2 U237 ( .A(n374), .B(n288), .Z(n284) );
  GTECH_NAND2 U238 ( .A(a[6]), .B(b[6]), .Z(n288) );
  GTECH_OAI21 U239 ( .A(a[6]), .B(b[6]), .C(n292), .Z(n374) );
  GTECH_OR_NOT U240 ( .A(n375), .B(n376), .Z(n292) );
  GTECH_OAI21 U241 ( .A(a[5]), .B(b[5]), .C(n299), .Z(n376) );
  GTECH_OR_NOT U242 ( .A(a[4]), .B(n301), .Z(n299) );
  GTECH_NOT U243 ( .A(b[4]), .Z(n301) );
  GTECH_NOT U244 ( .A(n294), .Z(n375) );
  GTECH_NAND2 U245 ( .A(a[5]), .B(b[5]), .Z(n294) );
  GTECH_XNOR2 U246 ( .A(a[4]), .B(b[4]), .Z(n302) );
  GTECH_AOI21 U247 ( .A(n356), .B(a[11]), .C(n377), .Z(n368) );
  GTECH_OA21 U248 ( .A(a[11]), .B(n356), .C(b[11]), .Z(n377) );
  GTECH_OAI21 U249 ( .A(n352), .B(n362), .C(n354), .Z(n356) );
  GTECH_NAND2 U250 ( .A(b[10]), .B(a[10]), .Z(n354) );
  GTECH_NOT U251 ( .A(n378), .Z(n362) );
  GTECH_AOI21 U252 ( .A(n276), .B(n275), .C(n361), .Z(n378) );
  GTECH_NOR2 U253 ( .A(b[9]), .B(a[9]), .Z(n361) );
  GTECH_NOR2 U254 ( .A(a[8]), .B(b[8]), .Z(n275) );
  GTECH_NAND2 U255 ( .A(b[9]), .B(a[9]), .Z(n276) );
  GTECH_NOR2 U256 ( .A(a[10]), .B(b[10]), .Z(n352) );
endmodule

