
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392;

  GTECH_MUX2 U139 ( .A(n278), .B(n279), .S(n280), .Z(sum[9]) );
  GTECH_XOR2 U140 ( .A(n281), .B(n282), .Z(n279) );
  GTECH_XOR2 U141 ( .A(n283), .B(n282), .Z(n278) );
  GTECH_AOI21 U142 ( .A(a[9]), .B(b[9]), .C(n284), .Z(n282) );
  GTECH_XOR2 U143 ( .A(n285), .B(n286), .Z(sum[8]) );
  GTECH_MUX2 U144 ( .A(n287), .B(n288), .S(n289), .Z(sum[7]) );
  GTECH_XNOR2 U145 ( .A(n290), .B(n291), .Z(n288) );
  GTECH_XOR2 U146 ( .A(n290), .B(n292), .Z(n287) );
  GTECH_AND_NOT U147 ( .A(n293), .B(n294), .Z(n292) );
  GTECH_OAI21 U148 ( .A(b[6]), .B(a[6]), .C(n295), .Z(n293) );
  GTECH_XNOR2 U149 ( .A(a[7]), .B(b[7]), .Z(n290) );
  GTECH_OAI21 U150 ( .A(n296), .B(n297), .C(n298), .Z(sum[6]) );
  GTECH_MUX2 U151 ( .A(n299), .B(n300), .S(b[6]), .Z(n298) );
  GTECH_OR_NOT U152 ( .A(a[6]), .B(n296), .Z(n300) );
  GTECH_XNOR2 U153 ( .A(a[6]), .B(n301), .Z(n299) );
  GTECH_NOT U154 ( .A(n294), .Z(n297) );
  GTECH_NOT U155 ( .A(n301), .Z(n296) );
  GTECH_AO21 U156 ( .A(n302), .B(n289), .C(n295), .Z(n301) );
  GTECH_OAI22 U157 ( .A(n303), .B(n304), .C(n305), .D(n306), .Z(n295) );
  GTECH_MUX2 U158 ( .A(n307), .B(n308), .S(n309), .Z(sum[5]) );
  GTECH_AOI21 U159 ( .A(a[5]), .B(b[5]), .C(n305), .Z(n309) );
  GTECH_OAI21 U160 ( .A(a[4]), .B(n289), .C(n310), .Z(n308) );
  GTECH_AO21 U161 ( .A(n289), .B(a[4]), .C(b[4]), .Z(n310) );
  GTECH_OAI21 U162 ( .A(n311), .B(n312), .C(n306), .Z(n307) );
  GTECH_NOT U163 ( .A(n313), .Z(n306) );
  GTECH_NOT U164 ( .A(n289), .Z(n312) );
  GTECH_XNOR2 U165 ( .A(n289), .B(n314), .Z(sum[4]) );
  GTECH_MUX2 U166 ( .A(n315), .B(n316), .S(n317), .Z(sum[3]) );
  GTECH_XOR2 U167 ( .A(n318), .B(n319), .Z(n316) );
  GTECH_AND2 U168 ( .A(n320), .B(n321), .Z(n319) );
  GTECH_AO21 U169 ( .A(n322), .B(n323), .C(n324), .Z(n321) );
  GTECH_XNOR2 U170 ( .A(n318), .B(n325), .Z(n315) );
  GTECH_XNOR2 U171 ( .A(a[3]), .B(b[3]), .Z(n318) );
  GTECH_MUX2 U172 ( .A(n326), .B(n327), .S(cin), .Z(sum[2]) );
  GTECH_MUX2 U173 ( .A(n328), .B(n329), .S(n330), .Z(n327) );
  GTECH_MUX2 U174 ( .A(n328), .B(n329), .S(n324), .Z(n326) );
  GTECH_OA21 U175 ( .A(n331), .B(n332), .C(n333), .Z(n324) );
  GTECH_XNOR2 U176 ( .A(a[2]), .B(n322), .Z(n329) );
  GTECH_OAI21 U177 ( .A(b[2]), .B(a[2]), .C(n320), .Z(n328) );
  GTECH_MUX2 U178 ( .A(n334), .B(n335), .S(n336), .Z(sum[1]) );
  GTECH_NOR2 U179 ( .A(n337), .B(n331), .Z(n336) );
  GTECH_AO21 U180 ( .A(n317), .B(n332), .C(n338), .Z(n335) );
  GTECH_OAI21 U181 ( .A(n338), .B(n317), .C(n332), .Z(n334) );
  GTECH_MUX2 U182 ( .A(n339), .B(n340), .S(n341), .Z(sum[15]) );
  GTECH_XNOR2 U183 ( .A(n342), .B(n343), .Z(n340) );
  GTECH_XOR2 U184 ( .A(n342), .B(n344), .Z(n339) );
  GTECH_AOI21 U185 ( .A(n345), .B(n346), .C(n347), .Z(n344) );
  GTECH_XNOR2 U186 ( .A(a[15]), .B(b[15]), .Z(n342) );
  GTECH_MUX2 U187 ( .A(n348), .B(n349), .S(n341), .Z(sum[14]) );
  GTECH_XNOR2 U188 ( .A(n350), .B(n351), .Z(n349) );
  GTECH_XNOR2 U189 ( .A(n350), .B(n346), .Z(n348) );
  GTECH_OA21 U190 ( .A(n352), .B(n353), .C(n354), .Z(n346) );
  GTECH_OR_NOT U191 ( .A(n347), .B(n345), .Z(n350) );
  GTECH_MUX2 U192 ( .A(n355), .B(n356), .S(n341), .Z(sum[13]) );
  GTECH_XNOR2 U193 ( .A(n357), .B(n358), .Z(n356) );
  GTECH_XNOR2 U194 ( .A(n353), .B(n357), .Z(n355) );
  GTECH_OAI21 U195 ( .A(a[13]), .B(b[13]), .C(n359), .Z(n357) );
  GTECH_NOT U196 ( .A(n352), .Z(n359) );
  GTECH_OAI21 U197 ( .A(n360), .B(n361), .C(n362), .Z(sum[12]) );
  GTECH_AND_NOT U198 ( .A(n358), .B(n353), .Z(n360) );
  GTECH_MUX2 U199 ( .A(n363), .B(n364), .S(n286), .Z(sum[11]) );
  GTECH_XNOR2 U200 ( .A(n365), .B(n366), .Z(n364) );
  GTECH_XOR2 U201 ( .A(n365), .B(n367), .Z(n363) );
  GTECH_AND_NOT U202 ( .A(n368), .B(n369), .Z(n367) );
  GTECH_OAI21 U203 ( .A(b[10]), .B(a[10]), .C(n370), .Z(n368) );
  GTECH_XNOR2 U204 ( .A(a[11]), .B(b[11]), .Z(n365) );
  GTECH_OAI21 U205 ( .A(n371), .B(n372), .C(n373), .Z(sum[10]) );
  GTECH_MUX2 U206 ( .A(n374), .B(n375), .S(b[10]), .Z(n373) );
  GTECH_OR_NOT U207 ( .A(a[10]), .B(n371), .Z(n375) );
  GTECH_XNOR2 U208 ( .A(a[10]), .B(n376), .Z(n374) );
  GTECH_NOT U209 ( .A(n369), .Z(n372) );
  GTECH_NOT U210 ( .A(n376), .Z(n371) );
  GTECH_AO21 U211 ( .A(n377), .B(n286), .C(n370), .Z(n376) );
  GTECH_AO22 U212 ( .A(a[9]), .B(b[9]), .C(n378), .D(n281), .Z(n370) );
  GTECH_NOT U213 ( .A(n280), .Z(n286) );
  GTECH_XNOR2 U214 ( .A(n317), .B(n379), .Z(sum[0]) );
  GTECH_OAI21 U215 ( .A(n380), .B(n361), .C(n362), .Z(cout) );
  GTECH_NAND3 U216 ( .A(n381), .B(n358), .C(n361), .Z(n362) );
  GTECH_NOT U217 ( .A(n353), .Z(n381) );
  GTECH_AND2 U218 ( .A(b[12]), .B(a[12]), .Z(n353) );
  GTECH_NOT U219 ( .A(n341), .Z(n361) );
  GTECH_MUX2 U220 ( .A(n382), .B(n285), .S(n280), .Z(n341) );
  GTECH_MUX2 U221 ( .A(n314), .B(n383), .S(n289), .Z(n280) );
  GTECH_MUX2 U222 ( .A(n384), .B(n379), .S(n317), .Z(n289) );
  GTECH_NOT U223 ( .A(cin), .Z(n317) );
  GTECH_AND_NOT U224 ( .A(n332), .B(n338), .Z(n379) );
  GTECH_OR_NOT U225 ( .A(n385), .B(b[0]), .Z(n332) );
  GTECH_OA21 U226 ( .A(a[3]), .B(n325), .C(n386), .Z(n384) );
  GTECH_AO21 U227 ( .A(n325), .B(a[3]), .C(b[3]), .Z(n386) );
  GTECH_OAI21 U228 ( .A(n330), .B(n387), .C(n320), .Z(n325) );
  GTECH_OR_NOT U229 ( .A(n323), .B(b[2]), .Z(n320) );
  GTECH_NOT U230 ( .A(a[2]), .Z(n323) );
  GTECH_AND_NOT U231 ( .A(n322), .B(a[2]), .Z(n387) );
  GTECH_NOT U232 ( .A(b[2]), .Z(n322) );
  GTECH_OA21 U233 ( .A(n331), .B(n338), .C(n333), .Z(n330) );
  GTECH_NOT U234 ( .A(n337), .Z(n333) );
  GTECH_AND2 U235 ( .A(a[1]), .B(b[1]), .Z(n337) );
  GTECH_AND_NOT U236 ( .A(n385), .B(b[0]), .Z(n338) );
  GTECH_NOT U237 ( .A(a[0]), .Z(n385) );
  GTECH_NOR2 U238 ( .A(a[1]), .B(b[1]), .Z(n331) );
  GTECH_AOI21 U239 ( .A(n291), .B(a[7]), .C(n388), .Z(n383) );
  GTECH_OA21 U240 ( .A(a[7]), .B(n291), .C(b[7]), .Z(n388) );
  GTECH_AO21 U241 ( .A(n302), .B(n389), .C(n294), .Z(n291) );
  GTECH_AND2 U242 ( .A(b[6]), .B(a[6]), .Z(n294) );
  GTECH_OR2 U243 ( .A(b[6]), .B(a[6]), .Z(n389) );
  GTECH_OAI22 U244 ( .A(n303), .B(n304), .C(n311), .D(n305), .Z(n302) );
  GTECH_AND_NOT U245 ( .A(n303), .B(b[5]), .Z(n305) );
  GTECH_NOT U246 ( .A(b[5]), .Z(n304) );
  GTECH_NOT U247 ( .A(a[5]), .Z(n303) );
  GTECH_OR2 U248 ( .A(n311), .B(n313), .Z(n314) );
  GTECH_AND2 U249 ( .A(a[4]), .B(b[4]), .Z(n313) );
  GTECH_NOR2 U250 ( .A(a[4]), .B(b[4]), .Z(n311) );
  GTECH_AND_NOT U251 ( .A(n283), .B(n281), .Z(n285) );
  GTECH_AND2 U252 ( .A(b[8]), .B(a[8]), .Z(n281) );
  GTECH_OA21 U253 ( .A(a[11]), .B(n366), .C(n390), .Z(n382) );
  GTECH_AO21 U254 ( .A(n366), .B(a[11]), .C(b[11]), .Z(n390) );
  GTECH_AO21 U255 ( .A(n377), .B(n391), .C(n369), .Z(n366) );
  GTECH_AND2 U256 ( .A(b[10]), .B(a[10]), .Z(n369) );
  GTECH_OR2 U257 ( .A(b[10]), .B(a[10]), .Z(n391) );
  GTECH_AO22 U258 ( .A(a[9]), .B(b[9]), .C(n283), .D(n378), .Z(n377) );
  GTECH_NOT U259 ( .A(n284), .Z(n378) );
  GTECH_NOR2 U260 ( .A(a[9]), .B(b[9]), .Z(n284) );
  GTECH_OR2 U261 ( .A(a[8]), .B(b[8]), .Z(n283) );
  GTECH_AOI21 U262 ( .A(n343), .B(a[15]), .C(n392), .Z(n380) );
  GTECH_OA21 U263 ( .A(a[15]), .B(n343), .C(b[15]), .Z(n392) );
  GTECH_AO21 U264 ( .A(n345), .B(n351), .C(n347), .Z(n343) );
  GTECH_AND2 U265 ( .A(b[14]), .B(a[14]), .Z(n347) );
  GTECH_OA21 U266 ( .A(n352), .B(n358), .C(n354), .Z(n351) );
  GTECH_OR2 U267 ( .A(a[13]), .B(b[13]), .Z(n354) );
  GTECH_OR2 U268 ( .A(a[12]), .B(b[12]), .Z(n358) );
  GTECH_AND2 U269 ( .A(b[13]), .B(a[13]), .Z(n352) );
  GTECH_OR2 U270 ( .A(a[14]), .B(b[14]), .Z(n345) );
endmodule

