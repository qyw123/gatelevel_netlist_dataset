
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NAND2 U83 ( .A(n93), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI21 U86 ( .A(n98), .B(n99), .C(n100), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n101), .B(n102), .C(n103), .Z(n100) );
  GTECH_NOT U88 ( .A(n102), .Z(n98) );
  GTECH_NAND2 U89 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n104), .Z(n84) );
  GTECH_NAND2 U91 ( .A(n105), .B(n106), .Z(n104) );
  GTECH_XOR2 U92 ( .A(n106), .B(n105), .Z(N153) );
  GTECH_NOT U93 ( .A(n107), .Z(n105) );
  GTECH_XOR3 U94 ( .A(n108), .B(n93), .C(n95), .Z(n107) );
  GTECH_XOR3 U95 ( .A(n101), .B(n103), .C(n102), .Z(n95) );
  GTECH_OAI21 U96 ( .A(n109), .B(n110), .C(n111), .Z(n102) );
  GTECH_OAI21 U97 ( .A(n112), .B(n113), .C(n114), .Z(n111) );
  GTECH_NOT U98 ( .A(n113), .Z(n109) );
  GTECH_NOT U99 ( .A(n115), .Z(n103) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n115) );
  GTECH_NOT U101 ( .A(n99), .Z(n101) );
  GTECH_NAND2 U102 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U103 ( .A(n116), .B(n117), .C(n118), .COUT(n93) );
  GTECH_NOT U104 ( .A(n119), .Z(n118) );
  GTECH_XOR2 U105 ( .A(n120), .B(n121), .Z(n117) );
  GTECH_AND2 U106 ( .A(I_a[7]), .B(I_b[5]), .Z(n121) );
  GTECH_NOT U107 ( .A(n122), .Z(n120) );
  GTECH_NOT U108 ( .A(n94), .Z(n108) );
  GTECH_NAND2 U109 ( .A(I_a[7]), .B(n122), .Z(n94) );
  GTECH_NOT U110 ( .A(n123), .Z(n106) );
  GTECH_NAND2 U111 ( .A(n124), .B(n125), .Z(n123) );
  GTECH_NOT U112 ( .A(n126), .Z(n125) );
  GTECH_XOR2 U113 ( .A(n126), .B(n127), .Z(N152) );
  GTECH_NOT U114 ( .A(n124), .Z(n127) );
  GTECH_XNOR4 U115 ( .A(n128), .B(n119), .C(n122), .D(n116), .Z(n124) );
  GTECH_ADD_ABC U116 ( .A(n129), .B(n130), .C(n131), .COUT(n116) );
  GTECH_NOT U117 ( .A(n132), .Z(n131) );
  GTECH_XOR3 U118 ( .A(n133), .B(n134), .C(n135), .Z(n130) );
  GTECH_OAI21 U119 ( .A(n135), .B(n136), .C(n137), .Z(n122) );
  GTECH_OAI21 U120 ( .A(n133), .B(n138), .C(n134), .Z(n137) );
  GTECH_NOT U121 ( .A(n138), .Z(n135) );
  GTECH_XOR3 U122 ( .A(n112), .B(n114), .C(n113), .Z(n119) );
  GTECH_OAI21 U123 ( .A(n139), .B(n140), .C(n141), .Z(n113) );
  GTECH_OAI21 U124 ( .A(n142), .B(n143), .C(n144), .Z(n141) );
  GTECH_NOT U125 ( .A(n143), .Z(n139) );
  GTECH_NOT U126 ( .A(n145), .Z(n114) );
  GTECH_NAND2 U127 ( .A(I_b[7]), .B(I_a[5]), .Z(n145) );
  GTECH_NOT U128 ( .A(n110), .Z(n112) );
  GTECH_NAND2 U129 ( .A(I_b[6]), .B(I_a[6]), .Z(n110) );
  GTECH_AND2 U130 ( .A(I_a[7]), .B(I_b[5]), .Z(n128) );
  GTECH_ADD_ABC U131 ( .A(n146), .B(n147), .C(n148), .COUT(n126) );
  GTECH_NOT U132 ( .A(n149), .Z(n148) );
  GTECH_AOI2N2 U133 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n147) );
  GTECH_OA21 U134 ( .A(n154), .B(n155), .C(n156), .Z(n146) );
  GTECH_XOR3 U135 ( .A(n157), .B(n149), .C(n158), .Z(N151) );
  GTECH_OA21 U136 ( .A(n154), .B(n155), .C(n156), .Z(n158) );
  GTECH_OAI21 U137 ( .A(n159), .B(n160), .C(n161), .Z(n156) );
  GTECH_XOR2 U138 ( .A(n162), .B(n129), .Z(n149) );
  GTECH_ADD_ABC U139 ( .A(n163), .B(n164), .C(n165), .COUT(n129) );
  GTECH_NOT U140 ( .A(n166), .Z(n165) );
  GTECH_XOR3 U141 ( .A(n167), .B(n168), .C(n169), .Z(n164) );
  GTECH_XNOR4 U142 ( .A(n134), .B(n138), .C(n132), .D(n133), .Z(n162) );
  GTECH_NOT U143 ( .A(n136), .Z(n133) );
  GTECH_NAND2 U144 ( .A(I_a[7]), .B(I_b[4]), .Z(n136) );
  GTECH_XOR3 U145 ( .A(n142), .B(n144), .C(n143), .Z(n132) );
  GTECH_OAI21 U146 ( .A(n170), .B(n171), .C(n172), .Z(n143) );
  GTECH_OAI21 U147 ( .A(n173), .B(n174), .C(n175), .Z(n172) );
  GTECH_NOT U148 ( .A(n174), .Z(n170) );
  GTECH_NOT U149 ( .A(n176), .Z(n144) );
  GTECH_NAND2 U150 ( .A(I_b[7]), .B(I_a[4]), .Z(n176) );
  GTECH_NOT U151 ( .A(n140), .Z(n142) );
  GTECH_NAND2 U152 ( .A(I_b[6]), .B(I_a[5]), .Z(n140) );
  GTECH_OAI21 U153 ( .A(n169), .B(n177), .C(n178), .Z(n138) );
  GTECH_OAI21 U154 ( .A(n167), .B(n179), .C(n168), .Z(n178) );
  GTECH_NOT U155 ( .A(n179), .Z(n169) );
  GTECH_NOT U156 ( .A(n180), .Z(n134) );
  GTECH_NAND2 U157 ( .A(I_a[6]), .B(I_b[5]), .Z(n180) );
  GTECH_AOI2N2 U158 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n157) );
  GTECH_NOT U159 ( .A(I_a[7]), .Z(n153) );
  GTECH_XOR3 U160 ( .A(n154), .B(n159), .C(n181), .Z(N150) );
  GTECH_NOT U161 ( .A(n161), .Z(n181) );
  GTECH_XOR2 U162 ( .A(n182), .B(n163), .Z(n161) );
  GTECH_ADD_ABC U163 ( .A(n183), .B(n184), .C(n185), .COUT(n163) );
  GTECH_NOT U164 ( .A(n186), .Z(n185) );
  GTECH_XOR3 U165 ( .A(n187), .B(n188), .C(n189), .Z(n184) );
  GTECH_XNOR4 U166 ( .A(n168), .B(n179), .C(n166), .D(n167), .Z(n182) );
  GTECH_NOT U167 ( .A(n177), .Z(n167) );
  GTECH_NAND2 U168 ( .A(I_a[6]), .B(I_b[4]), .Z(n177) );
  GTECH_XOR3 U169 ( .A(n173), .B(n175), .C(n174), .Z(n166) );
  GTECH_OAI21 U170 ( .A(n190), .B(n191), .C(n192), .Z(n174) );
  GTECH_OAI21 U171 ( .A(n193), .B(n194), .C(n195), .Z(n192) );
  GTECH_NOT U172 ( .A(n194), .Z(n190) );
  GTECH_NOT U173 ( .A(n196), .Z(n175) );
  GTECH_NAND2 U174 ( .A(I_b[7]), .B(I_a[3]), .Z(n196) );
  GTECH_NOT U175 ( .A(n171), .Z(n173) );
  GTECH_NAND2 U176 ( .A(I_b[6]), .B(I_a[4]), .Z(n171) );
  GTECH_OAI21 U177 ( .A(n189), .B(n197), .C(n198), .Z(n179) );
  GTECH_OAI21 U178 ( .A(n187), .B(n199), .C(n188), .Z(n198) );
  GTECH_NOT U179 ( .A(n199), .Z(n189) );
  GTECH_NOT U180 ( .A(n200), .Z(n168) );
  GTECH_NAND2 U181 ( .A(I_a[5]), .B(I_b[5]), .Z(n200) );
  GTECH_NOT U182 ( .A(n155), .Z(n159) );
  GTECH_XOR2 U183 ( .A(n150), .B(n201), .Z(n155) );
  GTECH_NOT U184 ( .A(n151), .Z(n201) );
  GTECH_OAI2N2 U185 ( .A(n202), .B(n203), .C(n204), .D(n205), .Z(n151) );
  GTECH_NAND2 U186 ( .A(n202), .B(n203), .Z(n205) );
  GTECH_XOR2 U187 ( .A(n206), .B(n152), .Z(n150) );
  GTECH_AND2 U188 ( .A(n207), .B(n208), .Z(n152) );
  GTECH_OR_NOT U189 ( .A(n209), .B(n210), .Z(n208) );
  GTECH_OAI21 U190 ( .A(n211), .B(n210), .C(n212), .Z(n207) );
  GTECH_NAND2 U191 ( .A(I_a[7]), .B(I_b[3]), .Z(n206) );
  GTECH_NOT U192 ( .A(n160), .Z(n154) );
  GTECH_OAI2N2 U193 ( .A(n213), .B(n214), .C(n215), .D(n216), .Z(n160) );
  GTECH_NAND2 U194 ( .A(n213), .B(n214), .Z(n216) );
  GTECH_XOR3 U195 ( .A(n213), .B(n217), .C(n218), .Z(N149) );
  GTECH_NOT U196 ( .A(n215), .Z(n218) );
  GTECH_XOR2 U197 ( .A(n219), .B(n183), .Z(n215) );
  GTECH_ADD_ABC U198 ( .A(n220), .B(n221), .C(n222), .COUT(n183) );
  GTECH_XOR3 U199 ( .A(n223), .B(n224), .C(n225), .Z(n221) );
  GTECH_OA21 U200 ( .A(n226), .B(n227), .C(n228), .Z(n220) );
  GTECH_XNOR4 U201 ( .A(n188), .B(n199), .C(n186), .D(n187), .Z(n219) );
  GTECH_NOT U202 ( .A(n197), .Z(n187) );
  GTECH_NAND2 U203 ( .A(I_a[5]), .B(I_b[4]), .Z(n197) );
  GTECH_XOR3 U204 ( .A(n193), .B(n195), .C(n194), .Z(n186) );
  GTECH_OAI21 U205 ( .A(n229), .B(n230), .C(n231), .Z(n194) );
  GTECH_NOT U206 ( .A(n232), .Z(n195) );
  GTECH_NAND2 U207 ( .A(I_b[7]), .B(I_a[2]), .Z(n232) );
  GTECH_NOT U208 ( .A(n191), .Z(n193) );
  GTECH_NAND2 U209 ( .A(I_b[6]), .B(I_a[3]), .Z(n191) );
  GTECH_OAI21 U210 ( .A(n225), .B(n233), .C(n234), .Z(n199) );
  GTECH_OAI21 U211 ( .A(n223), .B(n235), .C(n224), .Z(n234) );
  GTECH_NOT U212 ( .A(n235), .Z(n225) );
  GTECH_NOT U213 ( .A(n236), .Z(n188) );
  GTECH_NAND2 U214 ( .A(I_b[5]), .B(I_a[4]), .Z(n236) );
  GTECH_NOT U215 ( .A(n214), .Z(n217) );
  GTECH_XOR3 U216 ( .A(n237), .B(n202), .C(n204), .Z(n214) );
  GTECH_XOR3 U217 ( .A(n211), .B(n212), .C(n210), .Z(n204) );
  GTECH_OAI21 U218 ( .A(n238), .B(n239), .C(n240), .Z(n210) );
  GTECH_OAI21 U219 ( .A(n241), .B(n242), .C(n243), .Z(n240) );
  GTECH_NOT U220 ( .A(n242), .Z(n238) );
  GTECH_NOT U221 ( .A(n244), .Z(n212) );
  GTECH_NAND2 U222 ( .A(I_a[6]), .B(I_b[3]), .Z(n244) );
  GTECH_NOT U223 ( .A(n209), .Z(n211) );
  GTECH_NAND2 U224 ( .A(I_a[7]), .B(I_b[2]), .Z(n209) );
  GTECH_ADD_ABC U225 ( .A(n245), .B(n246), .C(n247), .COUT(n202) );
  GTECH_XOR2 U226 ( .A(n248), .B(n249), .Z(n246) );
  GTECH_AND2 U227 ( .A(I_a[7]), .B(I_b[1]), .Z(n249) );
  GTECH_NOT U228 ( .A(n203), .Z(n237) );
  GTECH_NAND2 U229 ( .A(I_a[7]), .B(n250), .Z(n203) );
  GTECH_ADD_ABC U230 ( .A(n251), .B(n252), .C(n253), .COUT(n213) );
  GTECH_XOR3 U231 ( .A(n245), .B(n254), .C(n247), .Z(n252) );
  GTECH_NOT U232 ( .A(n255), .Z(n247) );
  GTECH_XOR3 U233 ( .A(n256), .B(n253), .C(n251), .Z(N148) );
  GTECH_ADD_ABC U234 ( .A(n257), .B(n258), .C(n259), .COUT(n251) );
  GTECH_NOT U235 ( .A(n260), .Z(n259) );
  GTECH_XOR3 U236 ( .A(n261), .B(n262), .C(n263), .Z(n258) );
  GTECH_XOR2 U237 ( .A(n264), .B(n265), .Z(n253) );
  GTECH_OA21 U238 ( .A(n226), .B(n227), .C(n228), .Z(n265) );
  GTECH_OAI21 U239 ( .A(n266), .B(n267), .C(n268), .Z(n228) );
  GTECH_NOT U240 ( .A(n226), .Z(n267) );
  GTECH_XNOR4 U241 ( .A(n224), .B(n235), .C(n222), .D(n223), .Z(n264) );
  GTECH_NOT U242 ( .A(n233), .Z(n223) );
  GTECH_NAND2 U243 ( .A(I_b[4]), .B(I_a[4]), .Z(n233) );
  GTECH_XOR3 U244 ( .A(n269), .B(n270), .C(n231), .Z(n222) );
  GTECH_NAND3 U245 ( .A(I_b[6]), .B(I_a[1]), .C(n271), .Z(n231) );
  GTECH_NOT U246 ( .A(n230), .Z(n270) );
  GTECH_NAND2 U247 ( .A(I_b[7]), .B(I_a[1]), .Z(n230) );
  GTECH_NOT U248 ( .A(n229), .Z(n269) );
  GTECH_NAND2 U249 ( .A(I_b[6]), .B(I_a[2]), .Z(n229) );
  GTECH_OAI21 U250 ( .A(n272), .B(n273), .C(n274), .Z(n235) );
  GTECH_OAI21 U251 ( .A(n275), .B(n276), .C(n277), .Z(n274) );
  GTECH_NOT U252 ( .A(n276), .Z(n272) );
  GTECH_NOT U253 ( .A(n278), .Z(n224) );
  GTECH_NAND2 U254 ( .A(I_b[5]), .B(I_a[3]), .Z(n278) );
  GTECH_XOR3 U255 ( .A(n254), .B(n255), .C(n245), .Z(n256) );
  GTECH_ADD_ABC U256 ( .A(n261), .B(n279), .C(n263), .COUT(n245) );
  GTECH_NOT U257 ( .A(n280), .Z(n263) );
  GTECH_XOR3 U258 ( .A(n281), .B(n282), .C(n283), .Z(n279) );
  GTECH_XOR3 U259 ( .A(n241), .B(n243), .C(n242), .Z(n255) );
  GTECH_OAI21 U260 ( .A(n284), .B(n285), .C(n286), .Z(n242) );
  GTECH_OAI21 U261 ( .A(n287), .B(n288), .C(n289), .Z(n286) );
  GTECH_NOT U262 ( .A(n288), .Z(n284) );
  GTECH_NOT U263 ( .A(n290), .Z(n243) );
  GTECH_NAND2 U264 ( .A(I_a[5]), .B(I_b[3]), .Z(n290) );
  GTECH_NOT U265 ( .A(n239), .Z(n241) );
  GTECH_NAND2 U266 ( .A(I_a[6]), .B(I_b[2]), .Z(n239) );
  GTECH_XOR2 U267 ( .A(n291), .B(n248), .Z(n254) );
  GTECH_NOT U268 ( .A(n250), .Z(n248) );
  GTECH_OAI21 U269 ( .A(n283), .B(n292), .C(n293), .Z(n250) );
  GTECH_OAI21 U270 ( .A(n281), .B(n294), .C(n282), .Z(n293) );
  GTECH_NOT U271 ( .A(n294), .Z(n283) );
  GTECH_AND2 U272 ( .A(I_a[7]), .B(I_b[1]), .Z(n291) );
  GTECH_XOR2 U273 ( .A(n295), .B(n257), .Z(N147) );
  GTECH_ADD_ABC U274 ( .A(n296), .B(n297), .C(n298), .COUT(n257) );
  GTECH_XOR3 U275 ( .A(n299), .B(n300), .C(n301), .Z(n297) );
  GTECH_NOT U276 ( .A(n302), .Z(n300) );
  GTECH_OA21 U277 ( .A(n303), .B(n304), .C(n305), .Z(n296) );
  GTECH_XNOR4 U278 ( .A(n262), .B(n280), .C(n260), .D(n261), .Z(n295) );
  GTECH_ADD_ABC U279 ( .A(n299), .B(n306), .C(n301), .COUT(n261) );
  GTECH_NOT U280 ( .A(n307), .Z(n301) );
  GTECH_XOR3 U281 ( .A(n308), .B(n309), .C(n310), .Z(n306) );
  GTECH_XOR3 U282 ( .A(n268), .B(n227), .C(n226), .Z(n260) );
  GTECH_XOR2 U283 ( .A(n311), .B(n271), .Z(n226) );
  GTECH_NOT U284 ( .A(n312), .Z(n271) );
  GTECH_NAND2 U285 ( .A(I_b[7]), .B(I_a[0]), .Z(n312) );
  GTECH_NAND2 U286 ( .A(I_b[6]), .B(I_a[1]), .Z(n311) );
  GTECH_NOT U287 ( .A(n266), .Z(n227) );
  GTECH_XOR3 U288 ( .A(n275), .B(n277), .C(n276), .Z(n266) );
  GTECH_OAI21 U289 ( .A(n313), .B(n314), .C(n315), .Z(n276) );
  GTECH_NOT U290 ( .A(n316), .Z(n277) );
  GTECH_NAND2 U291 ( .A(I_b[5]), .B(I_a[2]), .Z(n316) );
  GTECH_NOT U292 ( .A(n273), .Z(n275) );
  GTECH_NAND2 U293 ( .A(I_b[4]), .B(I_a[3]), .Z(n273) );
  GTECH_NOT U294 ( .A(n317), .Z(n268) );
  GTECH_NAND3 U295 ( .A(I_a[0]), .B(n318), .C(I_b[6]), .Z(n317) );
  GTECH_NOT U296 ( .A(n319), .Z(n318) );
  GTECH_XOR3 U297 ( .A(n287), .B(n289), .C(n288), .Z(n280) );
  GTECH_OAI21 U298 ( .A(n320), .B(n321), .C(n322), .Z(n288) );
  GTECH_OAI21 U299 ( .A(n323), .B(n324), .C(n325), .Z(n322) );
  GTECH_NOT U300 ( .A(n324), .Z(n320) );
  GTECH_NOT U301 ( .A(n326), .Z(n289) );
  GTECH_NAND2 U302 ( .A(I_b[3]), .B(I_a[4]), .Z(n326) );
  GTECH_NOT U303 ( .A(n285), .Z(n287) );
  GTECH_NAND2 U304 ( .A(I_a[5]), .B(I_b[2]), .Z(n285) );
  GTECH_NOT U305 ( .A(n327), .Z(n262) );
  GTECH_XOR3 U306 ( .A(n281), .B(n282), .C(n294), .Z(n327) );
  GTECH_OAI21 U307 ( .A(n310), .B(n328), .C(n329), .Z(n294) );
  GTECH_OAI21 U308 ( .A(n308), .B(n330), .C(n309), .Z(n329) );
  GTECH_NOT U309 ( .A(n330), .Z(n310) );
  GTECH_NOT U310 ( .A(n331), .Z(n282) );
  GTECH_NAND2 U311 ( .A(I_a[6]), .B(I_b[1]), .Z(n331) );
  GTECH_NOT U312 ( .A(n292), .Z(n281) );
  GTECH_NAND2 U313 ( .A(I_a[7]), .B(I_b[0]), .Z(n292) );
  GTECH_XOR2 U314 ( .A(n332), .B(n333), .Z(N146) );
  GTECH_XNOR4 U315 ( .A(n307), .B(n299), .C(n302), .D(n298), .Z(n333) );
  GTECH_XOR2 U316 ( .A(n319), .B(n334), .Z(n298) );
  GTECH_AND2 U317 ( .A(I_b[6]), .B(I_a[0]), .Z(n334) );
  GTECH_XOR3 U318 ( .A(n335), .B(n336), .C(n315), .Z(n319) );
  GTECH_NAND3 U319 ( .A(I_b[4]), .B(I_a[1]), .C(n337), .Z(n315) );
  GTECH_NOT U320 ( .A(n314), .Z(n336) );
  GTECH_NAND2 U321 ( .A(I_b[5]), .B(I_a[1]), .Z(n314) );
  GTECH_NOT U322 ( .A(n313), .Z(n335) );
  GTECH_NAND2 U323 ( .A(I_b[4]), .B(I_a[2]), .Z(n313) );
  GTECH_XOR3 U324 ( .A(n308), .B(n309), .C(n330), .Z(n302) );
  GTECH_OAI21 U325 ( .A(n338), .B(n339), .C(n340), .Z(n330) );
  GTECH_OAI21 U326 ( .A(n341), .B(n342), .C(n343), .Z(n340) );
  GTECH_NOT U327 ( .A(n344), .Z(n309) );
  GTECH_NAND2 U328 ( .A(I_a[5]), .B(I_b[1]), .Z(n344) );
  GTECH_NOT U329 ( .A(n328), .Z(n308) );
  GTECH_NAND2 U330 ( .A(I_a[6]), .B(I_b[0]), .Z(n328) );
  GTECH_ADD_ABC U331 ( .A(n345), .B(n346), .C(n347), .COUT(n299) );
  GTECH_NOT U332 ( .A(n348), .Z(n347) );
  GTECH_XOR3 U333 ( .A(n341), .B(n343), .C(n338), .Z(n346) );
  GTECH_NOT U334 ( .A(n342), .Z(n338) );
  GTECH_XOR3 U335 ( .A(n323), .B(n325), .C(n324), .Z(n307) );
  GTECH_OAI21 U336 ( .A(n349), .B(n350), .C(n351), .Z(n324) );
  GTECH_OAI21 U337 ( .A(n352), .B(n353), .C(n354), .Z(n351) );
  GTECH_NOT U338 ( .A(n353), .Z(n349) );
  GTECH_NOT U339 ( .A(n355), .Z(n325) );
  GTECH_NAND2 U340 ( .A(I_b[3]), .B(I_a[3]), .Z(n355) );
  GTECH_NOT U341 ( .A(n321), .Z(n323) );
  GTECH_NAND2 U342 ( .A(I_b[2]), .B(I_a[4]), .Z(n321) );
  GTECH_OA21 U343 ( .A(n303), .B(n304), .C(n305), .Z(n332) );
  GTECH_OAI21 U344 ( .A(n356), .B(n357), .C(n358), .Z(n305) );
  GTECH_NOT U345 ( .A(n303), .Z(n357) );
  GTECH_XOR3 U346 ( .A(n358), .B(n304), .C(n303), .Z(N145) );
  GTECH_XOR2 U347 ( .A(n359), .B(n337), .Z(n303) );
  GTECH_NOT U348 ( .A(n360), .Z(n337) );
  GTECH_NAND2 U349 ( .A(I_b[5]), .B(I_a[0]), .Z(n360) );
  GTECH_NAND2 U350 ( .A(I_b[4]), .B(I_a[1]), .Z(n359) );
  GTECH_NOT U351 ( .A(n356), .Z(n304) );
  GTECH_XOR2 U352 ( .A(n361), .B(n345), .Z(n356) );
  GTECH_ADD_ABC U353 ( .A(n362), .B(n363), .C(n364), .COUT(n345) );
  GTECH_XOR3 U354 ( .A(n365), .B(n366), .C(n367), .Z(n363) );
  GTECH_OA21 U355 ( .A(n368), .B(n369), .C(n370), .Z(n362) );
  GTECH_XNOR4 U356 ( .A(n343), .B(n342), .C(n348), .D(n341), .Z(n361) );
  GTECH_NOT U357 ( .A(n339), .Z(n341) );
  GTECH_NAND2 U358 ( .A(I_a[5]), .B(I_b[0]), .Z(n339) );
  GTECH_XOR3 U359 ( .A(n352), .B(n354), .C(n353), .Z(n348) );
  GTECH_OAI21 U360 ( .A(n371), .B(n372), .C(n373), .Z(n353) );
  GTECH_NOT U361 ( .A(n374), .Z(n354) );
  GTECH_NAND2 U362 ( .A(I_b[3]), .B(I_a[2]), .Z(n374) );
  GTECH_NOT U363 ( .A(n350), .Z(n352) );
  GTECH_NAND2 U364 ( .A(I_b[2]), .B(I_a[3]), .Z(n350) );
  GTECH_OAI21 U365 ( .A(n367), .B(n375), .C(n376), .Z(n342) );
  GTECH_OAI21 U366 ( .A(n365), .B(n377), .C(n366), .Z(n376) );
  GTECH_NOT U367 ( .A(n375), .Z(n365) );
  GTECH_NOT U368 ( .A(n377), .Z(n367) );
  GTECH_NOT U369 ( .A(n378), .Z(n343) );
  GTECH_NAND2 U370 ( .A(I_a[4]), .B(I_b[1]), .Z(n378) );
  GTECH_NOT U371 ( .A(n379), .Z(n358) );
  GTECH_NAND3 U372 ( .A(I_a[0]), .B(n380), .C(I_b[4]), .Z(n379) );
  GTECH_XOR2 U373 ( .A(n381), .B(n380), .Z(N144) );
  GTECH_XOR2 U374 ( .A(n382), .B(n383), .Z(n380) );
  GTECH_XNOR4 U375 ( .A(n366), .B(n377), .C(n375), .D(n364), .Z(n383) );
  GTECH_XOR3 U376 ( .A(n384), .B(n385), .C(n373), .Z(n364) );
  GTECH_NAND3 U377 ( .A(I_b[2]), .B(I_a[1]), .C(n386), .Z(n373) );
  GTECH_NOT U378 ( .A(n372), .Z(n385) );
  GTECH_NAND2 U379 ( .A(I_b[3]), .B(I_a[1]), .Z(n372) );
  GTECH_NOT U380 ( .A(n371), .Z(n384) );
  GTECH_NAND2 U381 ( .A(I_b[2]), .B(I_a[2]), .Z(n371) );
  GTECH_NAND2 U382 ( .A(I_a[4]), .B(I_b[0]), .Z(n375) );
  GTECH_OAI21 U383 ( .A(n387), .B(n388), .C(n389), .Z(n377) );
  GTECH_OAI21 U384 ( .A(n390), .B(n391), .C(n392), .Z(n389) );
  GTECH_NOT U385 ( .A(n391), .Z(n387) );
  GTECH_NOT U386 ( .A(n393), .Z(n366) );
  GTECH_NAND2 U387 ( .A(I_a[3]), .B(I_b[1]), .Z(n393) );
  GTECH_OA21 U388 ( .A(n368), .B(n369), .C(n370), .Z(n382) );
  GTECH_OAI21 U389 ( .A(n394), .B(n395), .C(n396), .Z(n370) );
  GTECH_NOT U390 ( .A(n368), .Z(n395) );
  GTECH_AND2 U391 ( .A(I_b[4]), .B(I_a[0]), .Z(n381) );
  GTECH_XOR3 U392 ( .A(n396), .B(n369), .C(n368), .Z(N143) );
  GTECH_XOR2 U393 ( .A(n397), .B(n386), .Z(n368) );
  GTECH_NOT U394 ( .A(n398), .Z(n386) );
  GTECH_NAND2 U395 ( .A(I_b[3]), .B(I_a[0]), .Z(n398) );
  GTECH_NAND2 U396 ( .A(I_b[2]), .B(I_a[1]), .Z(n397) );
  GTECH_NOT U397 ( .A(n394), .Z(n369) );
  GTECH_XOR3 U398 ( .A(n390), .B(n392), .C(n391), .Z(n394) );
  GTECH_OAI21 U399 ( .A(n399), .B(n400), .C(n401), .Z(n391) );
  GTECH_NOT U400 ( .A(n402), .Z(n392) );
  GTECH_NAND2 U401 ( .A(I_b[1]), .B(I_a[2]), .Z(n402) );
  GTECH_NOT U402 ( .A(n388), .Z(n390) );
  GTECH_NAND2 U403 ( .A(I_b[0]), .B(I_a[3]), .Z(n388) );
  GTECH_NOT U404 ( .A(n403), .Z(n396) );
  GTECH_NAND3 U405 ( .A(I_a[0]), .B(n404), .C(I_b[2]), .Z(n403) );
  GTECH_XOR2 U406 ( .A(n405), .B(n404), .Z(N142) );
  GTECH_NOT U407 ( .A(n406), .Z(n404) );
  GTECH_XOR3 U408 ( .A(n407), .B(n408), .C(n401), .Z(n406) );
  GTECH_NAND3 U409 ( .A(n409), .B(I_b[0]), .C(I_a[1]), .Z(n401) );
  GTECH_NOT U410 ( .A(n399), .Z(n408) );
  GTECH_NAND2 U411 ( .A(I_a[1]), .B(I_b[1]), .Z(n399) );
  GTECH_NOT U412 ( .A(n400), .Z(n407) );
  GTECH_NAND2 U413 ( .A(I_b[0]), .B(I_a[2]), .Z(n400) );
  GTECH_AND2 U414 ( .A(I_b[2]), .B(I_a[0]), .Z(n405) );
  GTECH_XOR2 U415 ( .A(n409), .B(n410), .Z(N141) );
  GTECH_AND2 U416 ( .A(I_a[1]), .B(I_b[0]), .Z(n410) );
  GTECH_NOT U417 ( .A(n411), .Z(n409) );
  GTECH_NAND2 U418 ( .A(I_a[0]), .B(I_b[1]), .Z(n411) );
  GTECH_AND2 U419 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

