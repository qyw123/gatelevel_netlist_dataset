
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_AO21 U75 ( .A(n83), .B(n84), .C(n85), .Z(N155) );
  GTECH_OAI22 U76 ( .A(n86), .B(n87), .C(n88), .D(n89), .Z(n85) );
  GTECH_NOT U77 ( .A(n90), .Z(n89) );
  GTECH_XOR2 U78 ( .A(n83), .B(n84), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n84) );
  GTECH_XOR2 U80 ( .A(n90), .B(n88), .Z(n91) );
  GTECH_AOI2N2 U81 ( .A(n92), .B(n93), .C(n94), .D(n95), .Z(n88) );
  GTECH_NAND2 U82 ( .A(n94), .B(n95), .Z(n93) );
  GTECH_XOR2 U83 ( .A(n87), .B(n86), .Z(n90) );
  GTECH_OA21 U84 ( .A(n96), .B(n97), .C(n98), .Z(n86) );
  GTECH_AO21 U85 ( .A(n96), .B(n97), .C(n99), .Z(n98) );
  GTECH_NOT U86 ( .A(n100), .Z(n96) );
  GTECH_NAND2 U87 ( .A(I_b[7]), .B(I_a[7]), .Z(n87) );
  GTECH_NOT U88 ( .A(n101), .Z(n83) );
  GTECH_NAND2 U89 ( .A(n102), .B(n103), .Z(n101) );
  GTECH_XOR2 U90 ( .A(n103), .B(n102), .Z(N153) );
  GTECH_NOT U91 ( .A(n104), .Z(n102) );
  GTECH_XOR3 U92 ( .A(n105), .B(n94), .C(n92), .Z(n104) );
  GTECH_XOR3 U93 ( .A(n106), .B(n107), .C(n100), .Z(n92) );
  GTECH_OAI22 U94 ( .A(n108), .B(n109), .C(n110), .D(n111), .Z(n100) );
  GTECH_AND2 U95 ( .A(n108), .B(n109), .Z(n110) );
  GTECH_NOT U96 ( .A(n112), .Z(n108) );
  GTECH_NOT U97 ( .A(n99), .Z(n107) );
  GTECH_NAND2 U98 ( .A(I_b[7]), .B(I_a[6]), .Z(n99) );
  GTECH_NOT U99 ( .A(n97), .Z(n106) );
  GTECH_NAND2 U100 ( .A(I_a[7]), .B(I_b[6]), .Z(n97) );
  GTECH_ADD_ABC U101 ( .A(n113), .B(n114), .C(n115), .COUT(n94) );
  GTECH_NOT U102 ( .A(n116), .Z(n115) );
  GTECH_XOR2 U103 ( .A(n117), .B(n118), .Z(n114) );
  GTECH_AND2 U104 ( .A(I_a[7]), .B(I_b[5]), .Z(n118) );
  GTECH_NOT U105 ( .A(n95), .Z(n105) );
  GTECH_NAND2 U106 ( .A(I_a[7]), .B(n119), .Z(n95) );
  GTECH_NOT U107 ( .A(n120), .Z(n103) );
  GTECH_NAND2 U108 ( .A(n121), .B(n122), .Z(n120) );
  GTECH_NOT U109 ( .A(n123), .Z(n122) );
  GTECH_XOR2 U110 ( .A(n123), .B(n124), .Z(N152) );
  GTECH_NOT U111 ( .A(n121), .Z(n124) );
  GTECH_XOR4 U112 ( .A(n125), .B(n117), .C(n113), .D(n116), .Z(n121) );
  GTECH_XOR3 U113 ( .A(n126), .B(n127), .C(n112), .Z(n116) );
  GTECH_OAI22 U114 ( .A(n128), .B(n129), .C(n130), .D(n131), .Z(n112) );
  GTECH_AND2 U115 ( .A(n128), .B(n129), .Z(n130) );
  GTECH_NOT U116 ( .A(n132), .Z(n128) );
  GTECH_NOT U117 ( .A(n111), .Z(n127) );
  GTECH_NAND2 U118 ( .A(I_b[7]), .B(I_a[5]), .Z(n111) );
  GTECH_NOT U119 ( .A(n109), .Z(n126) );
  GTECH_NAND2 U120 ( .A(I_b[6]), .B(I_a[6]), .Z(n109) );
  GTECH_ADD_ABC U121 ( .A(n133), .B(n134), .C(n135), .COUT(n113) );
  GTECH_NOT U122 ( .A(n136), .Z(n135) );
  GTECH_XOR3 U123 ( .A(n137), .B(n138), .C(n139), .Z(n134) );
  GTECH_NOT U124 ( .A(n140), .Z(n137) );
  GTECH_NOT U125 ( .A(n119), .Z(n117) );
  GTECH_OAI22 U126 ( .A(n139), .B(n140), .C(n141), .D(n142), .Z(n119) );
  GTECH_AND2 U127 ( .A(n139), .B(n140), .Z(n141) );
  GTECH_NOT U128 ( .A(n143), .Z(n139) );
  GTECH_AND2 U129 ( .A(I_a[7]), .B(I_b[5]), .Z(n125) );
  GTECH_ADD_ABC U130 ( .A(n144), .B(n145), .C(n146), .COUT(n123) );
  GTECH_NOT U131 ( .A(n147), .Z(n146) );
  GTECH_OA22 U132 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n145) );
  GTECH_OA21 U133 ( .A(n152), .B(n153), .C(n154), .Z(n144) );
  GTECH_AO21 U134 ( .A(n152), .B(n153), .C(n155), .Z(n154) );
  GTECH_XOR3 U135 ( .A(n156), .B(n147), .C(n157), .Z(N151) );
  GTECH_OA21 U136 ( .A(n152), .B(n153), .C(n158), .Z(n157) );
  GTECH_AO21 U137 ( .A(n152), .B(n153), .C(n155), .Z(n158) );
  GTECH_XOR2 U138 ( .A(n159), .B(n133), .Z(n147) );
  GTECH_ADD_ABC U139 ( .A(n160), .B(n161), .C(n162), .COUT(n133) );
  GTECH_NOT U140 ( .A(n163), .Z(n162) );
  GTECH_XOR3 U141 ( .A(n164), .B(n165), .C(n166), .Z(n161) );
  GTECH_XOR4 U142 ( .A(n138), .B(n143), .C(n140), .D(n136), .Z(n159) );
  GTECH_XOR3 U143 ( .A(n167), .B(n168), .C(n132), .Z(n136) );
  GTECH_OAI22 U144 ( .A(n169), .B(n170), .C(n171), .D(n172), .Z(n132) );
  GTECH_AND2 U145 ( .A(n169), .B(n170), .Z(n171) );
  GTECH_NOT U146 ( .A(n173), .Z(n169) );
  GTECH_NOT U147 ( .A(n131), .Z(n168) );
  GTECH_NAND2 U148 ( .A(I_b[7]), .B(I_a[4]), .Z(n131) );
  GTECH_NOT U149 ( .A(n129), .Z(n167) );
  GTECH_NAND2 U150 ( .A(I_b[6]), .B(I_a[5]), .Z(n129) );
  GTECH_NAND2 U151 ( .A(I_a[7]), .B(I_b[4]), .Z(n140) );
  GTECH_OAI22 U152 ( .A(n166), .B(n174), .C(n175), .D(n176), .Z(n143) );
  GTECH_AND2 U153 ( .A(n166), .B(n174), .Z(n175) );
  GTECH_NOT U154 ( .A(n177), .Z(n166) );
  GTECH_NOT U155 ( .A(n142), .Z(n138) );
  GTECH_NAND2 U156 ( .A(I_a[6]), .B(I_b[5]), .Z(n142) );
  GTECH_OA22 U157 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(n156) );
  GTECH_NOT U158 ( .A(n178), .Z(n151) );
  GTECH_NOT U159 ( .A(I_a[7]), .Z(n149) );
  GTECH_XOR3 U160 ( .A(n152), .B(n179), .C(n155), .Z(N150) );
  GTECH_XOR2 U161 ( .A(n160), .B(n180), .Z(n155) );
  GTECH_XOR4 U162 ( .A(n165), .B(n177), .C(n163), .D(n164), .Z(n180) );
  GTECH_NOT U163 ( .A(n174), .Z(n164) );
  GTECH_NAND2 U164 ( .A(I_a[6]), .B(I_b[4]), .Z(n174) );
  GTECH_XOR3 U165 ( .A(n181), .B(n182), .C(n173), .Z(n163) );
  GTECH_OAI22 U166 ( .A(n183), .B(n184), .C(n185), .D(n186), .Z(n173) );
  GTECH_AND2 U167 ( .A(n183), .B(n184), .Z(n185) );
  GTECH_NOT U168 ( .A(n187), .Z(n183) );
  GTECH_NOT U169 ( .A(n172), .Z(n182) );
  GTECH_NAND2 U170 ( .A(I_b[7]), .B(I_a[3]), .Z(n172) );
  GTECH_NOT U171 ( .A(n170), .Z(n181) );
  GTECH_NAND2 U172 ( .A(I_b[6]), .B(I_a[4]), .Z(n170) );
  GTECH_OAI22 U173 ( .A(n188), .B(n189), .C(n190), .D(n191), .Z(n177) );
  GTECH_AND2 U174 ( .A(n188), .B(n189), .Z(n190) );
  GTECH_NOT U175 ( .A(n176), .Z(n165) );
  GTECH_NAND2 U176 ( .A(I_a[5]), .B(I_b[5]), .Z(n176) );
  GTECH_ADD_ABC U177 ( .A(n192), .B(n193), .C(n194), .COUT(n160) );
  GTECH_NOT U178 ( .A(n195), .Z(n194) );
  GTECH_XOR3 U179 ( .A(n196), .B(n197), .C(n188), .Z(n193) );
  GTECH_NOT U180 ( .A(n198), .Z(n188) );
  GTECH_NOT U181 ( .A(n153), .Z(n179) );
  GTECH_XOR2 U182 ( .A(n178), .B(n150), .Z(n153) );
  GTECH_AOI2N2 U183 ( .A(n199), .B(n200), .C(n201), .D(n202), .Z(n150) );
  GTECH_NAND2 U184 ( .A(n201), .B(n202), .Z(n200) );
  GTECH_XOR2 U185 ( .A(n203), .B(n148), .Z(n178) );
  GTECH_OA21 U186 ( .A(n204), .B(n205), .C(n206), .Z(n148) );
  GTECH_AO21 U187 ( .A(n204), .B(n205), .C(n207), .Z(n206) );
  GTECH_NOT U188 ( .A(n208), .Z(n204) );
  GTECH_NAND2 U189 ( .A(I_a[7]), .B(I_b[3]), .Z(n203) );
  GTECH_OA21 U190 ( .A(n209), .B(n210), .C(n211), .Z(n152) );
  GTECH_AO21 U191 ( .A(n209), .B(n210), .C(n212), .Z(n211) );
  GTECH_XOR3 U192 ( .A(n209), .B(n213), .C(n212), .Z(N149) );
  GTECH_XOR2 U193 ( .A(n192), .B(n214), .Z(n212) );
  GTECH_XOR4 U194 ( .A(n197), .B(n198), .C(n195), .D(n196), .Z(n214) );
  GTECH_NOT U195 ( .A(n189), .Z(n196) );
  GTECH_NAND2 U196 ( .A(I_a[5]), .B(I_b[4]), .Z(n189) );
  GTECH_XOR3 U197 ( .A(n215), .B(n216), .C(n187), .Z(n195) );
  GTECH_AO21 U198 ( .A(n217), .B(n218), .C(n219), .Z(n187) );
  GTECH_NOT U199 ( .A(n220), .Z(n219) );
  GTECH_NOT U200 ( .A(n186), .Z(n216) );
  GTECH_NAND2 U201 ( .A(I_b[7]), .B(I_a[2]), .Z(n186) );
  GTECH_NOT U202 ( .A(n184), .Z(n215) );
  GTECH_NAND2 U203 ( .A(I_b[6]), .B(I_a[3]), .Z(n184) );
  GTECH_OAI22 U204 ( .A(n221), .B(n222), .C(n223), .D(n224), .Z(n198) );
  GTECH_AND2 U205 ( .A(n221), .B(n222), .Z(n223) );
  GTECH_NOT U206 ( .A(n191), .Z(n197) );
  GTECH_NAND2 U207 ( .A(I_b[5]), .B(I_a[4]), .Z(n191) );
  GTECH_ADD_ABC U208 ( .A(n225), .B(n226), .C(n227), .COUT(n192) );
  GTECH_XOR3 U209 ( .A(n228), .B(n229), .C(n221), .Z(n226) );
  GTECH_NOT U210 ( .A(n230), .Z(n221) );
  GTECH_NOT U211 ( .A(n222), .Z(n228) );
  GTECH_OA21 U212 ( .A(n231), .B(n232), .C(n233), .Z(n225) );
  GTECH_AO21 U213 ( .A(n231), .B(n232), .C(n234), .Z(n233) );
  GTECH_NOT U214 ( .A(n210), .Z(n213) );
  GTECH_XOR3 U215 ( .A(n235), .B(n201), .C(n199), .Z(n210) );
  GTECH_XOR3 U216 ( .A(n236), .B(n237), .C(n208), .Z(n199) );
  GTECH_OAI22 U217 ( .A(n238), .B(n239), .C(n240), .D(n241), .Z(n208) );
  GTECH_AND2 U218 ( .A(n238), .B(n239), .Z(n240) );
  GTECH_NOT U219 ( .A(n242), .Z(n238) );
  GTECH_NOT U220 ( .A(n207), .Z(n237) );
  GTECH_NAND2 U221 ( .A(I_a[6]), .B(I_b[3]), .Z(n207) );
  GTECH_NOT U222 ( .A(n205), .Z(n236) );
  GTECH_NAND2 U223 ( .A(I_a[7]), .B(I_b[2]), .Z(n205) );
  GTECH_ADD_ABC U224 ( .A(n243), .B(n244), .C(n245), .COUT(n201) );
  GTECH_XOR2 U225 ( .A(n246), .B(n247), .Z(n244) );
  GTECH_AND2 U226 ( .A(I_a[7]), .B(I_b[1]), .Z(n247) );
  GTECH_NOT U227 ( .A(n202), .Z(n235) );
  GTECH_NAND2 U228 ( .A(I_a[7]), .B(n248), .Z(n202) );
  GTECH_ADD_ABC U229 ( .A(n249), .B(n250), .C(n251), .COUT(n209) );
  GTECH_XOR3 U230 ( .A(n243), .B(n252), .C(n245), .Z(n250) );
  GTECH_NOT U231 ( .A(n253), .Z(n245) );
  GTECH_XOR2 U232 ( .A(n249), .B(n254), .Z(N148) );
  GTECH_XOR4 U233 ( .A(n252), .B(n253), .C(n251), .D(n243), .Z(n254) );
  GTECH_ADD_ABC U234 ( .A(n255), .B(n256), .C(n257), .COUT(n243) );
  GTECH_XOR3 U235 ( .A(n258), .B(n259), .C(n260), .Z(n256) );
  GTECH_XOR2 U236 ( .A(n261), .B(n262), .Z(n251) );
  GTECH_OA21 U237 ( .A(n231), .B(n232), .C(n263), .Z(n262) );
  GTECH_AO21 U238 ( .A(n231), .B(n232), .C(n234), .Z(n263) );
  GTECH_XOR4 U239 ( .A(n229), .B(n230), .C(n222), .D(n227), .Z(n261) );
  GTECH_XOR3 U240 ( .A(n218), .B(n217), .C(n220), .Z(n227) );
  GTECH_NAND3 U241 ( .A(I_b[6]), .B(I_a[1]), .C(n264), .Z(n220) );
  GTECH_NOT U242 ( .A(n265), .Z(n217) );
  GTECH_NAND2 U243 ( .A(I_b[7]), .B(I_a[1]), .Z(n265) );
  GTECH_NOT U244 ( .A(n266), .Z(n218) );
  GTECH_NAND2 U245 ( .A(I_b[6]), .B(I_a[2]), .Z(n266) );
  GTECH_NAND2 U246 ( .A(I_b[4]), .B(I_a[4]), .Z(n222) );
  GTECH_OAI22 U247 ( .A(n267), .B(n268), .C(n269), .D(n270), .Z(n230) );
  GTECH_AND2 U248 ( .A(n267), .B(n268), .Z(n269) );
  GTECH_NOT U249 ( .A(n271), .Z(n267) );
  GTECH_NOT U250 ( .A(n224), .Z(n229) );
  GTECH_NAND2 U251 ( .A(I_b[5]), .B(I_a[3]), .Z(n224) );
  GTECH_XOR3 U252 ( .A(n272), .B(n273), .C(n242), .Z(n253) );
  GTECH_OAI22 U253 ( .A(n274), .B(n275), .C(n276), .D(n277), .Z(n242) );
  GTECH_AND2 U254 ( .A(n274), .B(n275), .Z(n276) );
  GTECH_NOT U255 ( .A(n278), .Z(n274) );
  GTECH_NOT U256 ( .A(n241), .Z(n273) );
  GTECH_NAND2 U257 ( .A(I_a[5]), .B(I_b[3]), .Z(n241) );
  GTECH_NOT U258 ( .A(n239), .Z(n272) );
  GTECH_NAND2 U259 ( .A(I_a[6]), .B(I_b[2]), .Z(n239) );
  GTECH_XOR2 U260 ( .A(n279), .B(n246), .Z(n252) );
  GTECH_NOT U261 ( .A(n248), .Z(n246) );
  GTECH_OAI22 U262 ( .A(n260), .B(n280), .C(n281), .D(n282), .Z(n248) );
  GTECH_AND2 U263 ( .A(n260), .B(n280), .Z(n281) );
  GTECH_NOT U264 ( .A(n283), .Z(n260) );
  GTECH_AND2 U265 ( .A(I_a[7]), .B(I_b[1]), .Z(n279) );
  GTECH_ADD_ABC U266 ( .A(n284), .B(n285), .C(n286), .COUT(n249) );
  GTECH_NOT U267 ( .A(n287), .Z(n286) );
  GTECH_XOR3 U268 ( .A(n255), .B(n288), .C(n257), .Z(n285) );
  GTECH_NOT U269 ( .A(n289), .Z(n257) );
  GTECH_NOT U270 ( .A(n290), .Z(n288) );
  GTECH_XOR2 U271 ( .A(n291), .B(n284), .Z(N147) );
  GTECH_ADD_ABC U272 ( .A(n292), .B(n293), .C(n294), .COUT(n284) );
  GTECH_XOR3 U273 ( .A(n295), .B(n296), .C(n297), .Z(n293) );
  GTECH_OA21 U274 ( .A(n298), .B(n299), .C(n300), .Z(n292) );
  GTECH_AO21 U275 ( .A(n298), .B(n299), .C(n301), .Z(n300) );
  GTECH_XOR4 U276 ( .A(n289), .B(n255), .C(n290), .D(n287), .Z(n291) );
  GTECH_XOR3 U277 ( .A(n302), .B(n232), .C(n231), .Z(n287) );
  GTECH_XOR2 U278 ( .A(n303), .B(n264), .Z(n231) );
  GTECH_NOT U279 ( .A(n304), .Z(n264) );
  GTECH_NAND2 U280 ( .A(I_b[7]), .B(I_a[0]), .Z(n304) );
  GTECH_NAND2 U281 ( .A(I_b[6]), .B(I_a[1]), .Z(n303) );
  GTECH_NOT U282 ( .A(n305), .Z(n232) );
  GTECH_XOR3 U283 ( .A(n306), .B(n307), .C(n271), .Z(n305) );
  GTECH_AO21 U284 ( .A(n308), .B(n309), .C(n310), .Z(n271) );
  GTECH_NOT U285 ( .A(n311), .Z(n310) );
  GTECH_NOT U286 ( .A(n270), .Z(n307) );
  GTECH_NAND2 U287 ( .A(I_b[5]), .B(I_a[2]), .Z(n270) );
  GTECH_NOT U288 ( .A(n268), .Z(n306) );
  GTECH_NAND2 U289 ( .A(I_b[4]), .B(I_a[3]), .Z(n268) );
  GTECH_NOT U290 ( .A(n234), .Z(n302) );
  GTECH_NAND3 U291 ( .A(I_a[0]), .B(n312), .C(I_b[6]), .Z(n234) );
  GTECH_NOT U292 ( .A(n313), .Z(n312) );
  GTECH_XOR3 U293 ( .A(n258), .B(n259), .C(n283), .Z(n290) );
  GTECH_OAI22 U294 ( .A(n314), .B(n315), .C(n316), .D(n317), .Z(n283) );
  GTECH_AND2 U295 ( .A(n314), .B(n315), .Z(n316) );
  GTECH_NOT U296 ( .A(n282), .Z(n259) );
  GTECH_NAND2 U297 ( .A(I_a[6]), .B(I_b[1]), .Z(n282) );
  GTECH_NOT U298 ( .A(n280), .Z(n258) );
  GTECH_NAND2 U299 ( .A(I_a[7]), .B(I_b[0]), .Z(n280) );
  GTECH_ADD_ABC U300 ( .A(n295), .B(n318), .C(n297), .COUT(n255) );
  GTECH_NOT U301 ( .A(n319), .Z(n297) );
  GTECH_XOR3 U302 ( .A(n320), .B(n321), .C(n314), .Z(n318) );
  GTECH_NOT U303 ( .A(n322), .Z(n314) );
  GTECH_XOR3 U304 ( .A(n323), .B(n324), .C(n278), .Z(n289) );
  GTECH_OAI22 U305 ( .A(n325), .B(n326), .C(n327), .D(n328), .Z(n278) );
  GTECH_AND2 U306 ( .A(n325), .B(n326), .Z(n327) );
  GTECH_NOT U307 ( .A(n329), .Z(n325) );
  GTECH_NOT U308 ( .A(n277), .Z(n324) );
  GTECH_NAND2 U309 ( .A(I_b[3]), .B(I_a[4]), .Z(n277) );
  GTECH_NOT U310 ( .A(n275), .Z(n323) );
  GTECH_NAND2 U311 ( .A(I_a[5]), .B(I_b[2]), .Z(n275) );
  GTECH_XOR2 U312 ( .A(n330), .B(n331), .Z(N146) );
  GTECH_XOR4 U313 ( .A(n296), .B(n319), .C(n294), .D(n295), .Z(n331) );
  GTECH_ADD_ABC U314 ( .A(n332), .B(n333), .C(n334), .COUT(n295) );
  GTECH_NOT U315 ( .A(n335), .Z(n334) );
  GTECH_XOR3 U316 ( .A(n336), .B(n337), .C(n338), .Z(n333) );
  GTECH_XOR2 U317 ( .A(n313), .B(n339), .Z(n294) );
  GTECH_AND2 U318 ( .A(I_b[6]), .B(I_a[0]), .Z(n339) );
  GTECH_XOR3 U319 ( .A(n309), .B(n308), .C(n311), .Z(n313) );
  GTECH_NAND3 U320 ( .A(I_b[4]), .B(I_a[1]), .C(n340), .Z(n311) );
  GTECH_NOT U321 ( .A(n341), .Z(n308) );
  GTECH_NAND2 U322 ( .A(I_b[5]), .B(I_a[1]), .Z(n341) );
  GTECH_NOT U323 ( .A(n342), .Z(n309) );
  GTECH_NAND2 U324 ( .A(I_b[4]), .B(I_a[2]), .Z(n342) );
  GTECH_XOR3 U325 ( .A(n343), .B(n344), .C(n329), .Z(n319) );
  GTECH_OAI22 U326 ( .A(n345), .B(n346), .C(n347), .D(n348), .Z(n329) );
  GTECH_AND2 U327 ( .A(n345), .B(n346), .Z(n347) );
  GTECH_NOT U328 ( .A(n349), .Z(n345) );
  GTECH_NOT U329 ( .A(n328), .Z(n344) );
  GTECH_NAND2 U330 ( .A(I_b[3]), .B(I_a[3]), .Z(n328) );
  GTECH_NOT U331 ( .A(n326), .Z(n343) );
  GTECH_NAND2 U332 ( .A(I_b[2]), .B(I_a[4]), .Z(n326) );
  GTECH_NOT U333 ( .A(n350), .Z(n296) );
  GTECH_XOR3 U334 ( .A(n320), .B(n321), .C(n322), .Z(n350) );
  GTECH_OAI22 U335 ( .A(n338), .B(n351), .C(n352), .D(n353), .Z(n322) );
  GTECH_AND2 U336 ( .A(n338), .B(n351), .Z(n352) );
  GTECH_NOT U337 ( .A(n354), .Z(n338) );
  GTECH_NOT U338 ( .A(n317), .Z(n321) );
  GTECH_NAND2 U339 ( .A(I_a[5]), .B(I_b[1]), .Z(n317) );
  GTECH_NOT U340 ( .A(n315), .Z(n320) );
  GTECH_NAND2 U341 ( .A(I_a[6]), .B(I_b[0]), .Z(n315) );
  GTECH_OA21 U342 ( .A(n298), .B(n299), .C(n355), .Z(n330) );
  GTECH_AO21 U343 ( .A(n298), .B(n299), .C(n301), .Z(n355) );
  GTECH_XOR3 U344 ( .A(n356), .B(n299), .C(n298), .Z(N145) );
  GTECH_XOR2 U345 ( .A(n357), .B(n340), .Z(n298) );
  GTECH_NOT U346 ( .A(n358), .Z(n340) );
  GTECH_NAND2 U347 ( .A(I_b[5]), .B(I_a[0]), .Z(n358) );
  GTECH_NAND2 U348 ( .A(I_b[4]), .B(I_a[1]), .Z(n357) );
  GTECH_XOR2 U349 ( .A(n332), .B(n359), .Z(n299) );
  GTECH_XOR4 U350 ( .A(n337), .B(n354), .C(n335), .D(n336), .Z(n359) );
  GTECH_NOT U351 ( .A(n351), .Z(n336) );
  GTECH_NAND2 U352 ( .A(I_a[5]), .B(I_b[0]), .Z(n351) );
  GTECH_XOR3 U353 ( .A(n360), .B(n361), .C(n349), .Z(n335) );
  GTECH_AO21 U354 ( .A(n362), .B(n363), .C(n364), .Z(n349) );
  GTECH_NOT U355 ( .A(n365), .Z(n364) );
  GTECH_NOT U356 ( .A(n348), .Z(n361) );
  GTECH_NAND2 U357 ( .A(I_b[3]), .B(I_a[2]), .Z(n348) );
  GTECH_NOT U358 ( .A(n346), .Z(n360) );
  GTECH_NAND2 U359 ( .A(I_b[2]), .B(I_a[3]), .Z(n346) );
  GTECH_OAI22 U360 ( .A(n366), .B(n367), .C(n368), .D(n369), .Z(n354) );
  GTECH_AND2 U361 ( .A(n366), .B(n367), .Z(n368) );
  GTECH_NOT U362 ( .A(n353), .Z(n337) );
  GTECH_NAND2 U363 ( .A(I_a[4]), .B(I_b[1]), .Z(n353) );
  GTECH_ADD_ABC U364 ( .A(n370), .B(n371), .C(n372), .COUT(n332) );
  GTECH_XOR3 U365 ( .A(n373), .B(n374), .C(n366), .Z(n371) );
  GTECH_NOT U366 ( .A(n375), .Z(n366) );
  GTECH_OA21 U367 ( .A(n376), .B(n377), .C(n378), .Z(n370) );
  GTECH_AO21 U368 ( .A(n376), .B(n377), .C(n379), .Z(n378) );
  GTECH_NOT U369 ( .A(n301), .Z(n356) );
  GTECH_NAND3 U370 ( .A(I_a[0]), .B(n380), .C(I_b[4]), .Z(n301) );
  GTECH_XOR2 U371 ( .A(n381), .B(n380), .Z(N144) );
  GTECH_XOR2 U372 ( .A(n382), .B(n383), .Z(n380) );
  GTECH_XOR4 U373 ( .A(n374), .B(n375), .C(n372), .D(n373), .Z(n383) );
  GTECH_NOT U374 ( .A(n367), .Z(n373) );
  GTECH_NAND2 U375 ( .A(I_a[4]), .B(I_b[0]), .Z(n367) );
  GTECH_XOR3 U376 ( .A(n363), .B(n362), .C(n365), .Z(n372) );
  GTECH_NAND3 U377 ( .A(I_b[2]), .B(I_a[1]), .C(n384), .Z(n365) );
  GTECH_NOT U378 ( .A(n385), .Z(n362) );
  GTECH_NAND2 U379 ( .A(I_b[3]), .B(I_a[1]), .Z(n385) );
  GTECH_NOT U380 ( .A(n386), .Z(n363) );
  GTECH_NAND2 U381 ( .A(I_b[2]), .B(I_a[2]), .Z(n386) );
  GTECH_OAI22 U382 ( .A(n387), .B(n388), .C(n389), .D(n390), .Z(n375) );
  GTECH_AND2 U383 ( .A(n387), .B(n388), .Z(n389) );
  GTECH_NOT U384 ( .A(n391), .Z(n387) );
  GTECH_NOT U385 ( .A(n369), .Z(n374) );
  GTECH_NAND2 U386 ( .A(I_a[3]), .B(I_b[1]), .Z(n369) );
  GTECH_OA21 U387 ( .A(n376), .B(n377), .C(n392), .Z(n382) );
  GTECH_AO21 U388 ( .A(n376), .B(n377), .C(n379), .Z(n392) );
  GTECH_AND2 U389 ( .A(I_b[4]), .B(I_a[0]), .Z(n381) );
  GTECH_XOR3 U390 ( .A(n393), .B(n377), .C(n376), .Z(N143) );
  GTECH_XOR2 U391 ( .A(n394), .B(n384), .Z(n376) );
  GTECH_NOT U392 ( .A(n395), .Z(n384) );
  GTECH_NAND2 U393 ( .A(I_b[3]), .B(I_a[0]), .Z(n395) );
  GTECH_NAND2 U394 ( .A(I_b[2]), .B(I_a[1]), .Z(n394) );
  GTECH_NOT U395 ( .A(n396), .Z(n377) );
  GTECH_XOR3 U396 ( .A(n397), .B(n398), .C(n391), .Z(n396) );
  GTECH_AO21 U397 ( .A(n399), .B(n400), .C(n401), .Z(n391) );
  GTECH_NOT U398 ( .A(n402), .Z(n401) );
  GTECH_NOT U399 ( .A(n390), .Z(n398) );
  GTECH_NAND2 U400 ( .A(I_b[1]), .B(I_a[2]), .Z(n390) );
  GTECH_NOT U401 ( .A(n388), .Z(n397) );
  GTECH_NAND2 U402 ( .A(I_b[0]), .B(I_a[3]), .Z(n388) );
  GTECH_NOT U403 ( .A(n379), .Z(n393) );
  GTECH_NAND3 U404 ( .A(I_a[0]), .B(n403), .C(I_b[2]), .Z(n379) );
  GTECH_XOR2 U405 ( .A(n404), .B(n403), .Z(N142) );
  GTECH_NOT U406 ( .A(n405), .Z(n403) );
  GTECH_XOR3 U407 ( .A(n399), .B(n400), .C(n402), .Z(n405) );
  GTECH_NAND3 U408 ( .A(n406), .B(I_b[0]), .C(I_a[1]), .Z(n402) );
  GTECH_NOT U409 ( .A(n407), .Z(n400) );
  GTECH_NAND2 U410 ( .A(I_a[1]), .B(I_b[1]), .Z(n407) );
  GTECH_NOT U411 ( .A(n408), .Z(n399) );
  GTECH_NAND2 U412 ( .A(I_b[0]), .B(I_a[2]), .Z(n408) );
  GTECH_AND2 U413 ( .A(I_b[2]), .B(I_a[0]), .Z(n404) );
  GTECH_XOR2 U414 ( .A(n406), .B(n409), .Z(N141) );
  GTECH_AND2 U415 ( .A(I_a[1]), .B(I_b[0]), .Z(n409) );
  GTECH_NOT U416 ( .A(n410), .Z(n406) );
  GTECH_NAND2 U417 ( .A(I_a[0]), .B(I_b[1]), .Z(n410) );
  GTECH_AND2 U418 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

