
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148;

  GTECH_XOR2 U94 ( .A(n75), .B(n76), .Z(sum[9]) );
  GTECH_XOR2 U95 ( .A(n77), .B(n78), .Z(sum[8]) );
  GTECH_XNOR2 U96 ( .A(n79), .B(n80), .Z(sum[7]) );
  GTECH_OA21 U97 ( .A(n81), .B(n82), .C(n83), .Z(n80) );
  GTECH_XNOR2 U98 ( .A(n84), .B(n81), .Z(sum[6]) );
  GTECH_AOI21 U99 ( .A(n85), .B(n86), .C(n87), .Z(n81) );
  GTECH_XOR2 U100 ( .A(n86), .B(n85), .Z(sum[5]) );
  GTECH_OAI21 U101 ( .A(n88), .B(n89), .C(n90), .Z(n85) );
  GTECH_XNOR2 U102 ( .A(n91), .B(n88), .Z(sum[4]) );
  GTECH_XNOR2 U103 ( .A(n92), .B(n93), .Z(sum[3]) );
  GTECH_OA21 U104 ( .A(n94), .B(n95), .C(n96), .Z(n93) );
  GTECH_NOT U105 ( .A(n97), .Z(n95) );
  GTECH_XNOR2 U106 ( .A(n94), .B(n97), .Z(sum[2]) );
  GTECH_AOI21 U107 ( .A(n98), .B(n99), .C(n100), .Z(n94) );
  GTECH_XOR2 U108 ( .A(n99), .B(n98), .Z(sum[1]) );
  GTECH_AO22 U109 ( .A(n101), .B(cin), .C(a[0]), .D(b[0]), .Z(n98) );
  GTECH_XNOR2 U110 ( .A(n102), .B(n103), .Z(sum[15]) );
  GTECH_AOI21 U111 ( .A(n104), .B(n105), .C(n106), .Z(n103) );
  GTECH_XOR2 U112 ( .A(n104), .B(n105), .Z(sum[14]) );
  GTECH_NOT U113 ( .A(n107), .Z(n104) );
  GTECH_AOI21 U114 ( .A(n108), .B(n109), .C(n110), .Z(n107) );
  GTECH_XOR2 U115 ( .A(n109), .B(n108), .Z(sum[13]) );
  GTECH_AO22 U116 ( .A(a[12]), .B(b[12]), .C(cout), .D(n111), .Z(n108) );
  GTECH_XOR2 U117 ( .A(n111), .B(cout), .Z(sum[12]) );
  GTECH_XNOR2 U118 ( .A(n112), .B(n113), .Z(sum[11]) );
  GTECH_AOI21 U119 ( .A(n114), .B(n115), .C(n116), .Z(n113) );
  GTECH_XOR2 U120 ( .A(n114), .B(n115), .Z(sum[10]) );
  GTECH_NOT U121 ( .A(n117), .Z(n114) );
  GTECH_AOI21 U122 ( .A(n76), .B(n75), .C(n118), .Z(n117) );
  GTECH_AO22 U123 ( .A(a[8]), .B(b[8]), .C(n78), .D(n77), .Z(n76) );
  GTECH_XOR2 U124 ( .A(cin), .B(n101), .Z(sum[0]) );
  GTECH_OAI21 U125 ( .A(n119), .B(n120), .C(n121), .Z(cout) );
  GTECH_NOT U126 ( .A(n78), .Z(n119) );
  GTECH_OAI21 U127 ( .A(n88), .B(n122), .C(n123), .Z(n78) );
  GTECH_AND2 U128 ( .A(n124), .B(n125), .Z(n88) );
  GTECH_NAND4 U129 ( .A(n126), .B(n97), .C(cin), .D(n127), .Z(n124) );
  GTECH_AND3 U130 ( .A(n92), .B(n99), .C(n101), .Z(n127) );
  GTECH_AND4 U131 ( .A(n128), .B(n126), .C(n129), .D(n130), .Z(Pm) );
  GTECH_AND4 U132 ( .A(n97), .B(n101), .C(n92), .D(n99), .Z(n130) );
  GTECH_XOR2 U133 ( .A(a[0]), .B(b[0]), .Z(n101) );
  GTECH_OAI21 U134 ( .A(n131), .B(n120), .C(n121), .Z(Gm) );
  GTECH_AOI21 U135 ( .A(b[15]), .B(a[15]), .C(n132), .Z(n121) );
  GTECH_OA21 U136 ( .A(n133), .B(n106), .C(n102), .Z(n132) );
  GTECH_NOT U137 ( .A(n134), .Z(n106) );
  GTECH_OA21 U138 ( .A(n135), .B(n110), .C(n105), .Z(n133) );
  GTECH_AND2 U139 ( .A(b[13]), .B(a[13]), .Z(n110) );
  GTECH_AND3 U140 ( .A(a[12]), .B(n109), .C(b[12]), .Z(n135) );
  GTECH_NOT U141 ( .A(n129), .Z(n120) );
  GTECH_AND4 U142 ( .A(n105), .B(n111), .C(n102), .D(n109), .Z(n129) );
  GTECH_XOR2 U143 ( .A(a[13]), .B(b[13]), .Z(n109) );
  GTECH_XOR2 U144 ( .A(a[15]), .B(b[15]), .Z(n102) );
  GTECH_XOR2 U145 ( .A(a[12]), .B(b[12]), .Z(n111) );
  GTECH_OA21 U146 ( .A(a[14]), .B(b[14]), .C(n134), .Z(n105) );
  GTECH_NAND2 U147 ( .A(a[14]), .B(b[14]), .Z(n134) );
  GTECH_OA21 U148 ( .A(n125), .B(n122), .C(n123), .Z(n131) );
  GTECH_AOI21 U149 ( .A(b[11]), .B(a[11]), .C(n136), .Z(n123) );
  GTECH_OA21 U150 ( .A(n137), .B(n116), .C(n112), .Z(n136) );
  GTECH_NOT U151 ( .A(n138), .Z(n116) );
  GTECH_OA21 U152 ( .A(n139), .B(n118), .C(n115), .Z(n137) );
  GTECH_AND2 U153 ( .A(a[9]), .B(b[9]), .Z(n118) );
  GTECH_AND3 U154 ( .A(a[8]), .B(n75), .C(b[8]), .Z(n139) );
  GTECH_NOT U155 ( .A(n128), .Z(n122) );
  GTECH_AND4 U156 ( .A(n115), .B(n77), .C(n112), .D(n75), .Z(n128) );
  GTECH_XOR2 U157 ( .A(a[9]), .B(b[9]), .Z(n75) );
  GTECH_XOR2 U158 ( .A(a[11]), .B(b[11]), .Z(n112) );
  GTECH_XOR2 U159 ( .A(a[8]), .B(b[8]), .Z(n77) );
  GTECH_OA21 U160 ( .A(a[10]), .B(b[10]), .C(n138), .Z(n115) );
  GTECH_NAND2 U161 ( .A(a[10]), .B(b[10]), .Z(n138) );
  GTECH_AOI222 U162 ( .A(n126), .B(n140), .C(b[7]), .D(a[7]), .E(n79), .F(n141), .Z(n125) );
  GTECH_OAI21 U163 ( .A(n142), .B(n82), .C(n83), .Z(n141) );
  GTECH_AOI21 U164 ( .A(n86), .B(n143), .C(n87), .Z(n142) );
  GTECH_AND2 U165 ( .A(b[5]), .B(a[5]), .Z(n87) );
  GTECH_NOT U166 ( .A(n90), .Z(n143) );
  GTECH_NOT U167 ( .A(n144), .Z(n140) );
  GTECH_AOI21 U168 ( .A(b[3]), .B(a[3]), .C(n145), .Z(n144) );
  GTECH_OA21 U169 ( .A(n146), .B(n147), .C(n92), .Z(n145) );
  GTECH_XOR2 U170 ( .A(a[3]), .B(b[3]), .Z(n92) );
  GTECH_NOT U171 ( .A(n96), .Z(n147) );
  GTECH_OA21 U172 ( .A(n148), .B(n100), .C(n97), .Z(n146) );
  GTECH_OA21 U173 ( .A(a[2]), .B(b[2]), .C(n96), .Z(n97) );
  GTECH_NAND2 U174 ( .A(a[2]), .B(b[2]), .Z(n96) );
  GTECH_AND2 U175 ( .A(a[1]), .B(b[1]), .Z(n100) );
  GTECH_AND3 U176 ( .A(a[0]), .B(n99), .C(b[0]), .Z(n148) );
  GTECH_XOR2 U177 ( .A(a[1]), .B(b[1]), .Z(n99) );
  GTECH_AND4 U178 ( .A(n91), .B(n84), .C(n86), .D(n79), .Z(n126) );
  GTECH_XOR2 U179 ( .A(a[7]), .B(b[7]), .Z(n79) );
  GTECH_XOR2 U180 ( .A(a[5]), .B(b[5]), .Z(n86) );
  GTECH_NOT U181 ( .A(n82), .Z(n84) );
  GTECH_OAI21 U182 ( .A(b[6]), .B(a[6]), .C(n83), .Z(n82) );
  GTECH_NAND2 U183 ( .A(a[6]), .B(b[6]), .Z(n83) );
  GTECH_NOT U184 ( .A(n89), .Z(n91) );
  GTECH_OAI21 U185 ( .A(b[4]), .B(a[4]), .C(n90), .Z(n89) );
  GTECH_NAND2 U186 ( .A(a[4]), .B(b[4]), .Z(n90) );
endmodule

