
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389;

  GTECH_MUX2 U142 ( .A(n281), .B(n282), .S(n283), .Z(sum[9]) );
  GTECH_XOR2 U143 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_XOR2 U144 ( .A(n285), .B(n286), .Z(n281) );
  GTECH_AOI21 U145 ( .A(a[9]), .B(b[9]), .C(n287), .Z(n285) );
  GTECH_NOT U146 ( .A(n288), .Z(n287) );
  GTECH_XOR2 U147 ( .A(n283), .B(n289), .Z(sum[8]) );
  GTECH_MUX2 U148 ( .A(n290), .B(n291), .S(n292), .Z(sum[7]) );
  GTECH_XOR2 U149 ( .A(n293), .B(n294), .Z(n291) );
  GTECH_XNOR2 U150 ( .A(n293), .B(n295), .Z(n290) );
  GTECH_AND2 U151 ( .A(n296), .B(n297), .Z(n295) );
  GTECH_AO21 U152 ( .A(n298), .B(n299), .C(n300), .Z(n296) );
  GTECH_XOR2 U153 ( .A(a[7]), .B(b[7]), .Z(n293) );
  GTECH_OAI21 U154 ( .A(n301), .B(n297), .C(n302), .Z(sum[6]) );
  GTECH_MUX2 U155 ( .A(n303), .B(n304), .S(n298), .Z(n302) );
  GTECH_XNOR2 U156 ( .A(n299), .B(n301), .Z(n304) );
  GTECH_NAND2 U157 ( .A(n301), .B(n299), .Z(n303) );
  GTECH_OA21 U158 ( .A(n305), .B(n306), .C(n300), .Z(n301) );
  GTECH_OAI21 U159 ( .A(n307), .B(n308), .C(n309), .Z(n300) );
  GTECH_MUX2 U160 ( .A(n310), .B(n311), .S(n312), .Z(sum[5]) );
  GTECH_AND_NOT U161 ( .A(n309), .B(n307), .Z(n312) );
  GTECH_OAI21 U162 ( .A(n308), .B(n292), .C(n313), .Z(n311) );
  GTECH_AO21 U163 ( .A(n313), .B(n292), .C(n308), .Z(n310) );
  GTECH_XNOR2 U164 ( .A(n314), .B(n305), .Z(sum[4]) );
  GTECH_MUX2 U165 ( .A(n315), .B(n316), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U166 ( .A(n317), .B(n318), .Z(n316) );
  GTECH_XNOR2 U167 ( .A(n317), .B(n319), .Z(n315) );
  GTECH_AND2 U168 ( .A(n320), .B(n321), .Z(n319) );
  GTECH_OAI21 U169 ( .A(b[2]), .B(a[2]), .C(n322), .Z(n320) );
  GTECH_XOR2 U170 ( .A(a[3]), .B(b[3]), .Z(n317) );
  GTECH_MUX2 U171 ( .A(n323), .B(n324), .S(n325), .Z(sum[2]) );
  GTECH_NOT U172 ( .A(cin), .Z(n325) );
  GTECH_MUX2 U173 ( .A(n326), .B(n327), .S(n322), .Z(n324) );
  GTECH_OA21 U174 ( .A(n328), .B(n329), .C(n330), .Z(n322) );
  GTECH_MUX2 U175 ( .A(n326), .B(n327), .S(n331), .Z(n323) );
  GTECH_OAI21 U176 ( .A(b[2]), .B(a[2]), .C(n321), .Z(n327) );
  GTECH_XOR2 U177 ( .A(a[2]), .B(b[2]), .Z(n326) );
  GTECH_MUX2 U178 ( .A(n332), .B(n333), .S(n334), .Z(sum[1]) );
  GTECH_AND_NOT U179 ( .A(n330), .B(n328), .Z(n334) );
  GTECH_OAI21 U180 ( .A(cin), .B(n329), .C(n335), .Z(n333) );
  GTECH_AO21 U181 ( .A(n335), .B(cin), .C(n329), .Z(n332) );
  GTECH_MUX2 U182 ( .A(n336), .B(n337), .S(n338), .Z(sum[15]) );
  GTECH_XOR2 U183 ( .A(n339), .B(n340), .Z(n337) );
  GTECH_OA21 U184 ( .A(n341), .B(n342), .C(n343), .Z(n340) );
  GTECH_XNOR2 U185 ( .A(n339), .B(n344), .Z(n336) );
  GTECH_XNOR2 U186 ( .A(a[15]), .B(b[15]), .Z(n339) );
  GTECH_MUX2 U187 ( .A(n345), .B(n346), .S(n347), .Z(sum[14]) );
  GTECH_OA21 U188 ( .A(n348), .B(n338), .C(n342), .Z(n347) );
  GTECH_OAI21 U189 ( .A(n349), .B(n350), .C(n351), .Z(n342) );
  GTECH_XOR2 U190 ( .A(b[14]), .B(a[14]), .Z(n346) );
  GTECH_NAND2 U191 ( .A(n343), .B(n352), .Z(n345) );
  GTECH_MUX2 U192 ( .A(n353), .B(n354), .S(n355), .Z(sum[13]) );
  GTECH_OA21 U193 ( .A(n350), .B(n356), .C(n357), .Z(n355) );
  GTECH_NAND2 U194 ( .A(n351), .B(n358), .Z(n354) );
  GTECH_XOR2 U195 ( .A(b[13]), .B(a[13]), .Z(n353) );
  GTECH_NAND2 U196 ( .A(n359), .B(n360), .Z(sum[12]) );
  GTECH_OAI21 U197 ( .A(n361), .B(n350), .C(n356), .Z(n359) );
  GTECH_MUX2 U198 ( .A(n362), .B(n363), .S(n283), .Z(sum[11]) );
  GTECH_XOR2 U199 ( .A(n364), .B(n365), .Z(n363) );
  GTECH_XNOR2 U200 ( .A(n364), .B(n366), .Z(n362) );
  GTECH_AND2 U201 ( .A(n367), .B(n368), .Z(n366) );
  GTECH_OAI21 U202 ( .A(b[10]), .B(a[10]), .C(n369), .Z(n367) );
  GTECH_XOR2 U203 ( .A(a[11]), .B(b[11]), .Z(n364) );
  GTECH_OAI21 U204 ( .A(n370), .B(n368), .C(n371), .Z(sum[10]) );
  GTECH_MUX2 U205 ( .A(n372), .B(n373), .S(b[10]), .Z(n371) );
  GTECH_OR2 U206 ( .A(n374), .B(a[10]), .Z(n373) );
  GTECH_XNOR2 U207 ( .A(a[10]), .B(n374), .Z(n372) );
  GTECH_NOT U208 ( .A(n370), .Z(n374) );
  GTECH_AOI21 U209 ( .A(n375), .B(n283), .C(n369), .Z(n370) );
  GTECH_AO22 U210 ( .A(a[9]), .B(b[9]), .C(n288), .D(n286), .Z(n369) );
  GTECH_XOR2 U211 ( .A(cin), .B(n376), .Z(sum[0]) );
  GTECH_OAI21 U212 ( .A(n377), .B(n338), .C(n360), .Z(cout) );
  GTECH_OR3 U213 ( .A(n350), .B(n361), .C(n356), .Z(n360) );
  GTECH_NOT U214 ( .A(n357), .Z(n361) );
  GTECH_AND2 U215 ( .A(b[12]), .B(a[12]), .Z(n350) );
  GTECH_NOT U216 ( .A(n356), .Z(n338) );
  GTECH_MUX2 U217 ( .A(n289), .B(n378), .S(n283), .Z(n356) );
  GTECH_MUX2 U218 ( .A(n314), .B(n379), .S(n292), .Z(n283) );
  GTECH_NOT U219 ( .A(n305), .Z(n292) );
  GTECH_MUX2 U220 ( .A(n380), .B(n381), .S(cin), .Z(n305) );
  GTECH_AOI21 U221 ( .A(n318), .B(a[3]), .C(n382), .Z(n381) );
  GTECH_OA21 U222 ( .A(a[3]), .B(n318), .C(b[3]), .Z(n382) );
  GTECH_NAND2 U223 ( .A(n383), .B(n321), .Z(n318) );
  GTECH_NAND2 U224 ( .A(b[2]), .B(a[2]), .Z(n321) );
  GTECH_OAI21 U225 ( .A(a[2]), .B(b[2]), .C(n331), .Z(n383) );
  GTECH_OA21 U226 ( .A(n328), .B(n335), .C(n330), .Z(n331) );
  GTECH_OR2 U227 ( .A(b[1]), .B(a[1]), .Z(n330) );
  GTECH_AND2 U228 ( .A(b[1]), .B(a[1]), .Z(n328) );
  GTECH_NOT U229 ( .A(n376), .Z(n380) );
  GTECH_AND_NOT U230 ( .A(n335), .B(n329), .Z(n376) );
  GTECH_AND2 U231 ( .A(a[0]), .B(b[0]), .Z(n329) );
  GTECH_OR2 U232 ( .A(b[0]), .B(a[0]), .Z(n335) );
  GTECH_OA21 U233 ( .A(a[7]), .B(n294), .C(n384), .Z(n379) );
  GTECH_AO21 U234 ( .A(n294), .B(a[7]), .C(b[7]), .Z(n384) );
  GTECH_NAND2 U235 ( .A(n385), .B(n297), .Z(n294) );
  GTECH_OR2 U236 ( .A(n299), .B(n298), .Z(n297) );
  GTECH_AO21 U237 ( .A(n299), .B(n298), .C(n306), .Z(n385) );
  GTECH_OAI21 U238 ( .A(n307), .B(n313), .C(n309), .Z(n306) );
  GTECH_OR2 U239 ( .A(a[5]), .B(b[5]), .Z(n309) );
  GTECH_AND2 U240 ( .A(a[5]), .B(b[5]), .Z(n307) );
  GTECH_NOT U241 ( .A(b[6]), .Z(n298) );
  GTECH_NOT U242 ( .A(a[6]), .Z(n299) );
  GTECH_AND_NOT U243 ( .A(n313), .B(n308), .Z(n314) );
  GTECH_AND2 U244 ( .A(b[4]), .B(a[4]), .Z(n308) );
  GTECH_OR2 U245 ( .A(a[4]), .B(b[4]), .Z(n313) );
  GTECH_OA21 U246 ( .A(a[11]), .B(n365), .C(n386), .Z(n378) );
  GTECH_AO21 U247 ( .A(n365), .B(a[11]), .C(b[11]), .Z(n386) );
  GTECH_NAND2 U248 ( .A(n387), .B(n368), .Z(n365) );
  GTECH_NAND2 U249 ( .A(b[10]), .B(a[10]), .Z(n368) );
  GTECH_OAI21 U250 ( .A(a[10]), .B(b[10]), .C(n375), .Z(n387) );
  GTECH_AO22 U251 ( .A(a[9]), .B(b[9]), .C(n288), .D(n284), .Z(n375) );
  GTECH_NOT U252 ( .A(n388), .Z(n284) );
  GTECH_OR2 U253 ( .A(b[9]), .B(a[9]), .Z(n288) );
  GTECH_NOR2 U254 ( .A(n388), .B(n286), .Z(n289) );
  GTECH_AND2 U255 ( .A(a[8]), .B(b[8]), .Z(n286) );
  GTECH_NOR2 U256 ( .A(b[8]), .B(a[8]), .Z(n388) );
  GTECH_AOI21 U257 ( .A(n344), .B(a[15]), .C(n389), .Z(n377) );
  GTECH_OA21 U258 ( .A(a[15]), .B(n344), .C(b[15]), .Z(n389) );
  GTECH_OAI21 U259 ( .A(n341), .B(n348), .C(n343), .Z(n344) );
  GTECH_NAND2 U260 ( .A(b[14]), .B(a[14]), .Z(n343) );
  GTECH_OAI21 U261 ( .A(n349), .B(n357), .C(n351), .Z(n348) );
  GTECH_OR2 U262 ( .A(a[13]), .B(b[13]), .Z(n351) );
  GTECH_OR2 U263 ( .A(b[12]), .B(a[12]), .Z(n357) );
  GTECH_NOT U264 ( .A(n358), .Z(n349) );
  GTECH_NAND2 U265 ( .A(b[13]), .B(a[13]), .Z(n358) );
  GTECH_NOT U266 ( .A(n352), .Z(n341) );
  GTECH_OR2 U267 ( .A(a[14]), .B(b[14]), .Z(n352) );
endmodule

