
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136;

  GTECH_XOR2 U88 ( .A(n69), .B(n70), .Z(sum[9]) );
  GTECH_XNOR2 U89 ( .A(n71), .B(n72), .Z(sum[8]) );
  GTECH_XNOR2 U90 ( .A(n73), .B(n74), .Z(sum[7]) );
  GTECH_OA21 U91 ( .A(n75), .B(n76), .C(n77), .Z(n74) );
  GTECH_XOR2 U92 ( .A(n76), .B(n75), .Z(sum[6]) );
  GTECH_OA21 U93 ( .A(n78), .B(n79), .C(n80), .Z(n75) );
  GTECH_XNOR2 U94 ( .A(n81), .B(n78), .Z(sum[5]) );
  GTECH_AOI21 U95 ( .A(n82), .B(n83), .C(n84), .Z(n78) );
  GTECH_XOR2 U96 ( .A(n82), .B(n83), .Z(sum[4]) );
  GTECH_XNOR2 U97 ( .A(n85), .B(n86), .Z(sum[3]) );
  GTECH_AOI21 U98 ( .A(n87), .B(n88), .C(n89), .Z(n86) );
  GTECH_XOR2 U99 ( .A(n87), .B(n88), .Z(sum[2]) );
  GTECH_AO22 U100 ( .A(b[1]), .B(a[1]), .C(n90), .D(n91), .Z(n87) );
  GTECH_XOR2 U101 ( .A(n91), .B(n90), .Z(sum[1]) );
  GTECH_AO22 U102 ( .A(n92), .B(cin), .C(a[0]), .D(b[0]), .Z(n90) );
  GTECH_XNOR2 U103 ( .A(n93), .B(n94), .Z(sum[15]) );
  GTECH_OAI21 U104 ( .A(n95), .B(n96), .C(n97), .Z(n93) );
  GTECH_XOR2 U105 ( .A(n96), .B(n95), .Z(sum[14]) );
  GTECH_OA21 U106 ( .A(n98), .B(n99), .C(n100), .Z(n95) );
  GTECH_XOR2 U107 ( .A(n99), .B(n98), .Z(sum[13]) );
  GTECH_OA21 U108 ( .A(n101), .B(n102), .C(n103), .Z(n98) );
  GTECH_NOT U109 ( .A(cout), .Z(n101) );
  GTECH_XNOR2 U110 ( .A(n102), .B(cout), .Z(sum[12]) );
  GTECH_XNOR2 U111 ( .A(n104), .B(n105), .Z(sum[11]) );
  GTECH_OAI21 U112 ( .A(n106), .B(n107), .C(n108), .Z(n104) );
  GTECH_XOR2 U113 ( .A(n107), .B(n106), .Z(sum[10]) );
  GTECH_OA21 U114 ( .A(n70), .B(n69), .C(n109), .Z(n106) );
  GTECH_OA21 U115 ( .A(n110), .B(n71), .C(n111), .Z(n70) );
  GTECH_XOR2 U116 ( .A(cin), .B(n92), .Z(sum[0]) );
  GTECH_AO21 U117 ( .A(n72), .B(n112), .C(n113), .Z(cout) );
  GTECH_NOT U118 ( .A(n110), .Z(n72) );
  GTECH_AOI21 U119 ( .A(n82), .B(n114), .C(n115), .Z(n110) );
  GTECH_AO21 U120 ( .A(n116), .B(cin), .C(n117), .Z(n82) );
  GTECH_AND3 U121 ( .A(n114), .B(n116), .C(n112), .Z(Pm) );
  GTECH_AND5 U122 ( .A(n85), .B(n91), .C(n92), .D(n118), .E(n88), .Z(n116) );
  GTECH_XOR2 U123 ( .A(a[0]), .B(b[0]), .Z(n92) );
  GTECH_AO21 U124 ( .A(n119), .B(n112), .C(n113), .Z(Gm) );
  GTECH_OAI21 U125 ( .A(n120), .B(n94), .C(n121), .Z(n113) );
  GTECH_OA21 U126 ( .A(n122), .B(n96), .C(n97), .Z(n120) );
  GTECH_OA21 U127 ( .A(n103), .B(n99), .C(n100), .Z(n122) );
  GTECH_NOR4 U128 ( .A(n102), .B(n94), .C(n96), .D(n99), .Z(n112) );
  GTECH_OAI21 U129 ( .A(b[13]), .B(a[13]), .C(n100), .Z(n99) );
  GTECH_NAND2 U130 ( .A(b[13]), .B(a[13]), .Z(n100) );
  GTECH_OAI21 U131 ( .A(b[14]), .B(a[14]), .C(n97), .Z(n96) );
  GTECH_NAND2 U132 ( .A(b[14]), .B(a[14]), .Z(n97) );
  GTECH_OAI21 U133 ( .A(b[15]), .B(a[15]), .C(n121), .Z(n94) );
  GTECH_NAND2 U134 ( .A(a[15]), .B(b[15]), .Z(n121) );
  GTECH_OAI21 U135 ( .A(b[12]), .B(a[12]), .C(n103), .Z(n102) );
  GTECH_NAND2 U136 ( .A(a[12]), .B(b[12]), .Z(n103) );
  GTECH_AO21 U137 ( .A(n117), .B(n114), .C(n115), .Z(n119) );
  GTECH_OAI21 U138 ( .A(n123), .B(n105), .C(n124), .Z(n115) );
  GTECH_OA21 U139 ( .A(n125), .B(n107), .C(n108), .Z(n123) );
  GTECH_OA21 U140 ( .A(n111), .B(n69), .C(n109), .Z(n125) );
  GTECH_NOR4 U141 ( .A(n71), .B(n105), .C(n107), .D(n69), .Z(n114) );
  GTECH_OAI21 U142 ( .A(b[9]), .B(a[9]), .C(n109), .Z(n69) );
  GTECH_NAND2 U143 ( .A(a[9]), .B(b[9]), .Z(n109) );
  GTECH_OAI21 U144 ( .A(b[10]), .B(a[10]), .C(n108), .Z(n107) );
  GTECH_NAND2 U145 ( .A(b[10]), .B(a[10]), .Z(n108) );
  GTECH_OAI21 U146 ( .A(b[11]), .B(a[11]), .C(n124), .Z(n105) );
  GTECH_NAND2 U147 ( .A(a[11]), .B(b[11]), .Z(n124) );
  GTECH_OAI21 U148 ( .A(b[8]), .B(a[8]), .C(n111), .Z(n71) );
  GTECH_NAND2 U149 ( .A(a[8]), .B(b[8]), .Z(n111) );
  GTECH_NOT U150 ( .A(n126), .Z(n117) );
  GTECH_AOI222 U151 ( .A(a[7]), .B(b[7]), .C(n118), .D(n127), .E(n73), .F(n128), .Z(n126) );
  GTECH_OAI21 U152 ( .A(n129), .B(n76), .C(n77), .Z(n128) );
  GTECH_NOT U153 ( .A(n130), .Z(n76) );
  GTECH_OA21 U154 ( .A(n79), .B(n131), .C(n80), .Z(n129) );
  GTECH_NAND2 U155 ( .A(a[5]), .B(b[5]), .Z(n80) );
  GTECH_OAI2N2 U156 ( .A(n132), .B(n133), .C(b[3]), .D(a[3]), .Z(n127) );
  GTECH_NOT U157 ( .A(n85), .Z(n133) );
  GTECH_XOR2 U158 ( .A(a[3]), .B(b[3]), .Z(n85) );
  GTECH_AOI21 U159 ( .A(n134), .B(n88), .C(n89), .Z(n132) );
  GTECH_OA21 U160 ( .A(a[2]), .B(b[2]), .C(n135), .Z(n88) );
  GTECH_NOT U161 ( .A(n89), .Z(n135) );
  GTECH_AND2 U162 ( .A(a[2]), .B(b[2]), .Z(n89) );
  GTECH_AO21 U163 ( .A(b[1]), .B(a[1]), .C(n136), .Z(n134) );
  GTECH_AND3 U164 ( .A(a[0]), .B(n91), .C(b[0]), .Z(n136) );
  GTECH_XOR2 U165 ( .A(a[1]), .B(b[1]), .Z(n91) );
  GTECH_AND4 U166 ( .A(n130), .B(n83), .C(n81), .D(n73), .Z(n118) );
  GTECH_XOR2 U167 ( .A(a[7]), .B(b[7]), .Z(n73) );
  GTECH_NOT U168 ( .A(n79), .Z(n81) );
  GTECH_XNOR2 U169 ( .A(a[5]), .B(b[5]), .Z(n79) );
  GTECH_OA21 U170 ( .A(b[4]), .B(a[4]), .C(n131), .Z(n83) );
  GTECH_NOT U171 ( .A(n84), .Z(n131) );
  GTECH_AND2 U172 ( .A(a[4]), .B(b[4]), .Z(n84) );
  GTECH_OA21 U173 ( .A(b[6]), .B(a[6]), .C(n77), .Z(n130) );
  GTECH_NAND2 U174 ( .A(b[6]), .B(a[6]), .Z(n77) );
endmodule

