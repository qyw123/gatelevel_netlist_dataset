
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141;

  GTECH_XOR2 U96 ( .A(n77), .B(n78), .Z(sum[9]) );
  GTECH_XOR2 U97 ( .A(n79), .B(n80), .Z(sum[8]) );
  GTECH_XNOR2 U98 ( .A(n81), .B(n82), .Z(sum[7]) );
  GTECH_OA21 U99 ( .A(n83), .B(n84), .C(n85), .Z(n82) );
  GTECH_XOR2 U100 ( .A(n84), .B(n83), .Z(sum[6]) );
  GTECH_OA21 U101 ( .A(n86), .B(n87), .C(n88), .Z(n83) );
  GTECH_XOR2 U102 ( .A(n87), .B(n86), .Z(sum[5]) );
  GTECH_OA21 U103 ( .A(n89), .B(n90), .C(n91), .Z(n86) );
  GTECH_XOR2 U104 ( .A(n90), .B(n89), .Z(sum[4]) );
  GTECH_XOR2 U105 ( .A(n92), .B(n93), .Z(sum[3]) );
  GTECH_OA21 U106 ( .A(n94), .B(n95), .C(n96), .Z(n93) );
  GTECH_XOR2 U107 ( .A(n95), .B(n94), .Z(sum[2]) );
  GTECH_OA21 U108 ( .A(n97), .B(n98), .C(n99), .Z(n94) );
  GTECH_XOR2 U109 ( .A(n98), .B(n97), .Z(sum[1]) );
  GTECH_AND2 U110 ( .A(n100), .B(n101), .Z(n97) );
  GTECH_XOR2 U111 ( .A(n102), .B(n103), .Z(sum[15]) );
  GTECH_OA21 U112 ( .A(n104), .B(n105), .C(n106), .Z(n103) );
  GTECH_XOR2 U113 ( .A(n105), .B(n104), .Z(sum[14]) );
  GTECH_OA21 U114 ( .A(n107), .B(n108), .C(n109), .Z(n104) );
  GTECH_XOR2 U115 ( .A(n108), .B(n107), .Z(sum[13]) );
  GTECH_OA21 U116 ( .A(n110), .B(n111), .C(n112), .Z(n107) );
  GTECH_XOR2 U117 ( .A(n110), .B(n111), .Z(sum[12]) );
  GTECH_NOT U118 ( .A(cout), .Z(n110) );
  GTECH_XNOR2 U119 ( .A(n113), .B(n114), .Z(sum[11]) );
  GTECH_OAI21 U120 ( .A(n115), .B(n116), .C(n117), .Z(n113) );
  GTECH_XOR2 U121 ( .A(n116), .B(n115), .Z(sum[10]) );
  GTECH_OA21 U122 ( .A(n78), .B(n77), .C(n118), .Z(n115) );
  GTECH_OA21 U123 ( .A(n80), .B(n79), .C(n119), .Z(n78) );
  GTECH_XNOR2 U124 ( .A(cin), .B(n120), .Z(sum[0]) );
  GTECH_OAI21 U125 ( .A(n80), .B(n121), .C(n122), .Z(cout) );
  GTECH_OA21 U126 ( .A(n89), .B(n123), .C(n124), .Z(n80) );
  GTECH_AND2 U127 ( .A(n125), .B(n126), .Z(n89) );
  GTECH_OR5 U128 ( .A(n98), .B(n92), .C(n95), .D(n101), .E(n127), .Z(n125) );
  GTECH_OR_NOT U129 ( .A(n120), .B(cin), .Z(n101) );
  GTECH_NOR4 U130 ( .A(n123), .B(n127), .C(n121), .D(n128), .Z(Pm) );
  GTECH_OR4 U131 ( .A(n95), .B(n98), .C(n120), .D(n92), .Z(n128) );
  GTECH_XNOR2 U132 ( .A(a[0]), .B(b[0]), .Z(n120) );
  GTECH_NOT U133 ( .A(n129), .Z(n127) );
  GTECH_OAI21 U134 ( .A(n130), .B(n121), .C(n122), .Z(Gm) );
  GTECH_AOI2N2 U135 ( .A(b[15]), .B(a[15]), .C(n131), .D(n102), .Z(n122) );
  GTECH_OA21 U136 ( .A(n132), .B(n105), .C(n106), .Z(n131) );
  GTECH_OA21 U137 ( .A(n112), .B(n108), .C(n109), .Z(n132) );
  GTECH_OR4 U138 ( .A(n111), .B(n105), .C(n108), .D(n102), .Z(n121) );
  GTECH_XNOR2 U139 ( .A(a[15]), .B(b[15]), .Z(n102) );
  GTECH_OAI21 U140 ( .A(b[13]), .B(a[13]), .C(n109), .Z(n108) );
  GTECH_NAND2 U141 ( .A(b[13]), .B(a[13]), .Z(n109) );
  GTECH_OAI21 U142 ( .A(b[14]), .B(a[14]), .C(n106), .Z(n105) );
  GTECH_NAND2 U143 ( .A(b[14]), .B(a[14]), .Z(n106) );
  GTECH_OAI21 U144 ( .A(b[12]), .B(a[12]), .C(n112), .Z(n111) );
  GTECH_NAND2 U145 ( .A(b[12]), .B(a[12]), .Z(n112) );
  GTECH_OA21 U146 ( .A(n126), .B(n123), .C(n124), .Z(n130) );
  GTECH_OA21 U147 ( .A(n133), .B(n114), .C(n134), .Z(n124) );
  GTECH_OA21 U148 ( .A(n135), .B(n116), .C(n117), .Z(n133) );
  GTECH_OA21 U149 ( .A(n119), .B(n77), .C(n118), .Z(n135) );
  GTECH_NAND2 U150 ( .A(b[8]), .B(a[8]), .Z(n119) );
  GTECH_OR4 U151 ( .A(n114), .B(n116), .C(n77), .D(n79), .Z(n123) );
  GTECH_XNOR2 U152 ( .A(a[8]), .B(b[8]), .Z(n79) );
  GTECH_OAI21 U153 ( .A(b[9]), .B(a[9]), .C(n118), .Z(n77) );
  GTECH_NAND2 U154 ( .A(b[9]), .B(a[9]), .Z(n118) );
  GTECH_OAI21 U155 ( .A(b[10]), .B(a[10]), .C(n117), .Z(n116) );
  GTECH_NAND2 U156 ( .A(b[10]), .B(a[10]), .Z(n117) );
  GTECH_OAI21 U157 ( .A(a[11]), .B(b[11]), .C(n134), .Z(n114) );
  GTECH_NAND2 U158 ( .A(b[11]), .B(a[11]), .Z(n134) );
  GTECH_AOI222 U159 ( .A(n129), .B(n136), .C(b[7]), .D(a[7]), .E(n81), .F(n137), .Z(n126) );
  GTECH_OAI21 U160 ( .A(n138), .B(n84), .C(n85), .Z(n137) );
  GTECH_OA21 U161 ( .A(n87), .B(n91), .C(n88), .Z(n138) );
  GTECH_OAI2N2 U162 ( .A(n139), .B(n92), .C(b[3]), .D(a[3]), .Z(n136) );
  GTECH_XNOR2 U163 ( .A(a[3]), .B(b[3]), .Z(n92) );
  GTECH_OA21 U164 ( .A(n140), .B(n95), .C(n96), .Z(n139) );
  GTECH_OAI21 U165 ( .A(b[2]), .B(a[2]), .C(n96), .Z(n95) );
  GTECH_NAND2 U166 ( .A(b[2]), .B(a[2]), .Z(n96) );
  GTECH_OA21 U167 ( .A(n100), .B(n98), .C(n99), .Z(n140) );
  GTECH_OAI21 U168 ( .A(b[1]), .B(a[1]), .C(n99), .Z(n98) );
  GTECH_NAND2 U169 ( .A(b[1]), .B(a[1]), .Z(n99) );
  GTECH_NAND2 U170 ( .A(b[0]), .B(a[0]), .Z(n100) );
  GTECH_NOR4 U171 ( .A(n90), .B(n84), .C(n87), .D(n141), .Z(n129) );
  GTECH_NOT U172 ( .A(n81), .Z(n141) );
  GTECH_XOR2 U173 ( .A(a[7]), .B(b[7]), .Z(n81) );
  GTECH_OAI21 U174 ( .A(b[5]), .B(a[5]), .C(n88), .Z(n87) );
  GTECH_NAND2 U175 ( .A(b[5]), .B(a[5]), .Z(n88) );
  GTECH_OAI21 U176 ( .A(b[6]), .B(a[6]), .C(n85), .Z(n84) );
  GTECH_NAND2 U177 ( .A(b[6]), .B(a[6]), .Z(n85) );
  GTECH_OAI21 U178 ( .A(b[4]), .B(a[4]), .C(n91), .Z(n90) );
  GTECH_NAND2 U179 ( .A(b[4]), .B(a[4]), .Z(n91) );
endmodule

