
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138;

  GTECH_XOR2 U90 ( .A(n71), .B(n72), .Z(sum[9]) );
  GTECH_XOR2 U91 ( .A(n73), .B(n74), .Z(sum[8]) );
  GTECH_XNOR2 U92 ( .A(n75), .B(n76), .Z(sum[7]) );
  GTECH_OAI21 U93 ( .A(n77), .B(n78), .C(n79), .Z(n75) );
  GTECH_XOR2 U94 ( .A(n78), .B(n77), .Z(sum[6]) );
  GTECH_OA21 U95 ( .A(n80), .B(n81), .C(n82), .Z(n77) );
  GTECH_XOR2 U96 ( .A(n81), .B(n80), .Z(sum[5]) );
  GTECH_OA21 U97 ( .A(n83), .B(n84), .C(n85), .Z(n80) );
  GTECH_XOR2 U98 ( .A(n84), .B(n83), .Z(sum[4]) );
  GTECH_XOR2 U99 ( .A(n86), .B(n87), .Z(sum[3]) );
  GTECH_OA21 U100 ( .A(n88), .B(n89), .C(n90), .Z(n87) );
  GTECH_XOR2 U101 ( .A(n88), .B(n89), .Z(sum[2]) );
  GTECH_AOI22 U102 ( .A(b[1]), .B(a[1]), .C(n91), .D(n92), .Z(n88) );
  GTECH_XOR2 U103 ( .A(n92), .B(n91), .Z(sum[1]) );
  GTECH_AO22 U104 ( .A(n93), .B(cin), .C(a[0]), .D(b[0]), .Z(n91) );
  GTECH_XNOR2 U105 ( .A(n94), .B(n95), .Z(sum[15]) );
  GTECH_OAI21 U106 ( .A(n96), .B(n97), .C(n98), .Z(n94) );
  GTECH_XOR2 U107 ( .A(n96), .B(n97), .Z(sum[14]) );
  GTECH_AOI2N2 U108 ( .A(b[13]), .B(a[13]), .C(n99), .D(n100), .Z(n96) );
  GTECH_XOR2 U109 ( .A(n100), .B(n99), .Z(sum[13]) );
  GTECH_OA21 U110 ( .A(n101), .B(n102), .C(n103), .Z(n99) );
  GTECH_XNOR2 U111 ( .A(n102), .B(cout), .Z(sum[12]) );
  GTECH_XNOR2 U112 ( .A(n104), .B(n105), .Z(sum[11]) );
  GTECH_OAI21 U113 ( .A(n106), .B(n107), .C(n108), .Z(n104) );
  GTECH_XOR2 U114 ( .A(n107), .B(n106), .Z(sum[10]) );
  GTECH_OA21 U115 ( .A(n72), .B(n71), .C(n109), .Z(n106) );
  GTECH_OA21 U116 ( .A(n74), .B(n73), .C(n110), .Z(n72) );
  GTECH_XOR2 U117 ( .A(cin), .B(n93), .Z(sum[0]) );
  GTECH_NOT U118 ( .A(n101), .Z(cout) );
  GTECH_OA21 U119 ( .A(n74), .B(n111), .C(n112), .Z(n101) );
  GTECH_OA21 U120 ( .A(n83), .B(n113), .C(n114), .Z(n74) );
  GTECH_AOI21 U121 ( .A(n115), .B(cin), .C(n116), .Z(n83) );
  GTECH_NOT U122 ( .A(n117), .Z(n115) );
  GTECH_NOR3 U123 ( .A(n111), .B(n117), .C(n113), .Z(Pm) );
  GTECH_OR5 U124 ( .A(n86), .B(n118), .C(n119), .D(n120), .E(n89), .Z(n117) );
  GTECH_NOT U125 ( .A(n93), .Z(n119) );
  GTECH_XOR2 U126 ( .A(a[0]), .B(b[0]), .Z(n93) );
  GTECH_OAI21 U127 ( .A(n121), .B(n111), .C(n112), .Z(Gm) );
  GTECH_OA21 U128 ( .A(n122), .B(n95), .C(n123), .Z(n112) );
  GTECH_OA21 U129 ( .A(n124), .B(n97), .C(n98), .Z(n122) );
  GTECH_AOI2N2 U130 ( .A(b[13]), .B(a[13]), .C(n100), .D(n103), .Z(n124) );
  GTECH_OR4 U131 ( .A(n102), .B(n95), .C(n97), .D(n100), .Z(n111) );
  GTECH_XNOR2 U132 ( .A(a[13]), .B(b[13]), .Z(n100) );
  GTECH_OAI21 U133 ( .A(b[14]), .B(a[14]), .C(n98), .Z(n97) );
  GTECH_NAND2 U134 ( .A(b[14]), .B(a[14]), .Z(n98) );
  GTECH_OAI21 U135 ( .A(b[15]), .B(a[15]), .C(n123), .Z(n95) );
  GTECH_NAND2 U136 ( .A(a[15]), .B(b[15]), .Z(n123) );
  GTECH_OAI21 U137 ( .A(b[12]), .B(a[12]), .C(n103), .Z(n102) );
  GTECH_NAND2 U138 ( .A(b[12]), .B(a[12]), .Z(n103) );
  GTECH_OA21 U139 ( .A(n125), .B(n113), .C(n114), .Z(n121) );
  GTECH_NOT U140 ( .A(n126), .Z(n114) );
  GTECH_OAI21 U141 ( .A(n127), .B(n105), .C(n128), .Z(n126) );
  GTECH_OA21 U142 ( .A(n129), .B(n107), .C(n108), .Z(n127) );
  GTECH_OA21 U143 ( .A(n110), .B(n71), .C(n109), .Z(n129) );
  GTECH_OR4 U144 ( .A(n73), .B(n105), .C(n107), .D(n71), .Z(n113) );
  GTECH_OAI21 U145 ( .A(b[9]), .B(a[9]), .C(n109), .Z(n71) );
  GTECH_NAND2 U146 ( .A(a[9]), .B(b[9]), .Z(n109) );
  GTECH_OAI21 U147 ( .A(b[10]), .B(a[10]), .C(n108), .Z(n107) );
  GTECH_NAND2 U148 ( .A(b[10]), .B(a[10]), .Z(n108) );
  GTECH_OAI21 U149 ( .A(b[11]), .B(a[11]), .C(n128), .Z(n105) );
  GTECH_NAND2 U150 ( .A(a[11]), .B(b[11]), .Z(n128) );
  GTECH_OAI21 U151 ( .A(b[8]), .B(a[8]), .C(n110), .Z(n73) );
  GTECH_NAND2 U152 ( .A(a[8]), .B(b[8]), .Z(n110) );
  GTECH_NOT U153 ( .A(n116), .Z(n125) );
  GTECH_OAI21 U154 ( .A(n130), .B(n120), .C(n131), .Z(n116) );
  GTECH_OA21 U155 ( .A(n132), .B(n76), .C(n133), .Z(n131) );
  GTECH_OA21 U156 ( .A(n134), .B(n78), .C(n79), .Z(n132) );
  GTECH_OA21 U157 ( .A(n81), .B(n85), .C(n82), .Z(n134) );
  GTECH_NAND2 U158 ( .A(a[5]), .B(b[5]), .Z(n82) );
  GTECH_OR4 U159 ( .A(n84), .B(n76), .C(n78), .D(n81), .Z(n120) );
  GTECH_XNOR2 U160 ( .A(a[5]), .B(b[5]), .Z(n81) );
  GTECH_OAI21 U161 ( .A(b[6]), .B(a[6]), .C(n79), .Z(n78) );
  GTECH_NAND2 U162 ( .A(b[6]), .B(a[6]), .Z(n79) );
  GTECH_OAI21 U163 ( .A(b[7]), .B(a[7]), .C(n133), .Z(n76) );
  GTECH_NAND2 U164 ( .A(a[7]), .B(b[7]), .Z(n133) );
  GTECH_OAI21 U165 ( .A(b[4]), .B(a[4]), .C(n85), .Z(n84) );
  GTECH_NAND2 U166 ( .A(a[4]), .B(b[4]), .Z(n85) );
  GTECH_AOI2N2 U167 ( .A(b[3]), .B(a[3]), .C(n135), .D(n86), .Z(n130) );
  GTECH_XNOR2 U168 ( .A(a[3]), .B(b[3]), .Z(n86) );
  GTECH_OA21 U169 ( .A(n136), .B(n89), .C(n90), .Z(n135) );
  GTECH_OAI21 U170 ( .A(a[2]), .B(b[2]), .C(n90), .Z(n89) );
  GTECH_NAND2 U171 ( .A(b[2]), .B(a[2]), .Z(n90) );
  GTECH_AOI21 U172 ( .A(b[1]), .B(a[1]), .C(n137), .Z(n136) );
  GTECH_NOT U173 ( .A(n138), .Z(n137) );
  GTECH_NAND3 U174 ( .A(a[0]), .B(n92), .C(b[0]), .Z(n138) );
  GTECH_NOT U175 ( .A(n118), .Z(n92) );
  GTECH_XNOR2 U176 ( .A(a[1]), .B(b[1]), .Z(n118) );
endmodule

