
module carry_select_adder8 ( a, b, cin, cout, sum );
  input [7:0] a;
  input [7:0] b;
  output [7:0] sum;
  input cin;
  output cout;
  wire   n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192;

  GTECH_MUX2 U72 ( .A(n141), .B(n142), .S(n143), .Z(sum[7]) );
  GTECH_XOR2 U73 ( .A(n144), .B(n145), .Z(n142) );
  GTECH_AO21 U74 ( .A(n146), .B(n147), .C(n148), .Z(n145) );
  GTECH_XOR2 U75 ( .A(n144), .B(n149), .Z(n141) );
  GTECH_XOR2 U76 ( .A(a[7]), .B(b[7]), .Z(n144) );
  GTECH_MUX2 U77 ( .A(n150), .B(n151), .S(n152), .Z(sum[6]) );
  GTECH_OA21 U78 ( .A(n153), .B(n143), .C(n154), .Z(n152) );
  GTECH_NOT U79 ( .A(n147), .Z(n154) );
  GTECH_OAI21 U80 ( .A(n155), .B(n156), .C(n157), .Z(n147) );
  GTECH_XOR2 U81 ( .A(b[6]), .B(a[6]), .Z(n151) );
  GTECH_OR_NOT U82 ( .A(n148), .B(n146), .Z(n150) );
  GTECH_MUX2 U83 ( .A(n158), .B(n159), .S(n160), .Z(sum[5]) );
  GTECH_OA21 U84 ( .A(n161), .B(n143), .C(n156), .Z(n160) );
  GTECH_XOR2 U85 ( .A(b[5]), .B(a[5]), .Z(n159) );
  GTECH_OR_NOT U86 ( .A(n155), .B(n157), .Z(n158) );
  GTECH_OAI21 U87 ( .A(n162), .B(n143), .C(n163), .Z(sum[4]) );
  GTECH_MUX2 U88 ( .A(n164), .B(n165), .S(n166), .Z(sum[3]) );
  GTECH_XOR2 U89 ( .A(n167), .B(n168), .Z(n165) );
  GTECH_OA21 U90 ( .A(a[2]), .B(n169), .C(n170), .Z(n167) );
  GTECH_AO21 U91 ( .A(n169), .B(a[2]), .C(b[2]), .Z(n170) );
  GTECH_XOR2 U92 ( .A(n168), .B(n171), .Z(n164) );
  GTECH_XOR2 U93 ( .A(a[3]), .B(b[3]), .Z(n168) );
  GTECH_MUX2 U94 ( .A(n172), .B(n173), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U95 ( .A(n174), .B(n175), .Z(n173) );
  GTECH_XOR2 U96 ( .A(n174), .B(n169), .Z(n172) );
  GTECH_NAND2 U97 ( .A(n176), .B(n177), .Z(n169) );
  GTECH_OR3 U98 ( .A(n178), .B(n179), .C(n180), .Z(n176) );
  GTECH_XOR2 U99 ( .A(a[2]), .B(b[2]), .Z(n174) );
  GTECH_XNOR3 U100 ( .A(b[1]), .B(n181), .C(n182), .Z(sum[1]) );
  GTECH_OAI2N2 U101 ( .A(n183), .B(n166), .C(b[0]), .D(a[0]), .Z(n182) );
  GTECH_XOR2 U102 ( .A(n166), .B(n184), .Z(sum[0]) );
  GTECH_OAI21 U103 ( .A(n185), .B(n143), .C(n163), .Z(cout) );
  GTECH_NAND2 U104 ( .A(n143), .B(n162), .Z(n163) );
  GTECH_AND_NOT U105 ( .A(n156), .B(n161), .Z(n162) );
  GTECH_NAND2 U106 ( .A(b[4]), .B(a[4]), .Z(n156) );
  GTECH_MUX2 U107 ( .A(n186), .B(n184), .S(n166), .Z(n143) );
  GTECH_NOT U108 ( .A(cin), .Z(n166) );
  GTECH_XOR2 U109 ( .A(a[0]), .B(n178), .Z(n184) );
  GTECH_NOT U110 ( .A(n187), .Z(n186) );
  GTECH_AO21 U111 ( .A(n171), .B(a[3]), .C(n188), .Z(n187) );
  GTECH_OA21 U112 ( .A(a[3]), .B(n171), .C(b[3]), .Z(n188) );
  GTECH_AO21 U113 ( .A(n175), .B(a[2]), .C(n189), .Z(n171) );
  GTECH_OA21 U114 ( .A(a[2]), .B(n175), .C(b[2]), .Z(n189) );
  GTECH_OAI21 U115 ( .A(n179), .B(n183), .C(n177), .Z(n175) );
  GTECH_NAND2 U116 ( .A(a[1]), .B(b[1]), .Z(n177) );
  GTECH_AND2 U117 ( .A(n180), .B(n178), .Z(n183) );
  GTECH_NOT U118 ( .A(b[0]), .Z(n178) );
  GTECH_NOT U119 ( .A(a[0]), .Z(n180) );
  GTECH_AND_NOT U120 ( .A(n181), .B(b[1]), .Z(n179) );
  GTECH_NOT U121 ( .A(a[1]), .Z(n181) );
  GTECH_NOT U122 ( .A(n190), .Z(n185) );
  GTECH_AO21 U123 ( .A(n149), .B(a[7]), .C(n191), .Z(n190) );
  GTECH_OA21 U124 ( .A(a[7]), .B(n149), .C(b[7]), .Z(n191) );
  GTECH_AO21 U125 ( .A(n146), .B(n192), .C(n148), .Z(n149) );
  GTECH_AND2 U126 ( .A(a[6]), .B(b[6]), .Z(n148) );
  GTECH_NOT U127 ( .A(n153), .Z(n192) );
  GTECH_OA21 U128 ( .A(n161), .B(n155), .C(n157), .Z(n153) );
  GTECH_NAND2 U129 ( .A(b[5]), .B(a[5]), .Z(n157) );
  GTECH_NOR2 U130 ( .A(a[5]), .B(b[5]), .Z(n155) );
  GTECH_NOR2 U131 ( .A(b[4]), .B(a[4]), .Z(n161) );
  GTECH_OR2 U132 ( .A(b[6]), .B(a[6]), .Z(n146) );
endmodule

