
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144;

  GTECH_XOR2 U92 ( .A(n73), .B(n74), .Z(sum[9]) );
  GTECH_XOR2 U93 ( .A(n75), .B(n76), .Z(sum[8]) );
  GTECH_XNOR2 U94 ( .A(n77), .B(n78), .Z(sum[7]) );
  GTECH_OA21 U95 ( .A(n79), .B(n80), .C(n81), .Z(n78) );
  GTECH_XNOR2 U96 ( .A(n79), .B(n82), .Z(sum[6]) );
  GTECH_AOI22 U97 ( .A(n83), .B(n84), .C(b[5]), .D(a[5]), .Z(n79) );
  GTECH_XOR2 U98 ( .A(n84), .B(n83), .Z(sum[5]) );
  GTECH_AO22 U99 ( .A(a[4]), .B(b[4]), .C(n85), .D(n86), .Z(n83) );
  GTECH_XOR2 U100 ( .A(n86), .B(n85), .Z(sum[4]) );
  GTECH_XOR2 U101 ( .A(n87), .B(n88), .Z(sum[3]) );
  GTECH_OA21 U102 ( .A(n89), .B(n90), .C(n91), .Z(n88) );
  GTECH_XNOR2 U103 ( .A(n89), .B(n92), .Z(sum[2]) );
  GTECH_AOI22 U104 ( .A(n93), .B(n94), .C(b[1]), .D(a[1]), .Z(n89) );
  GTECH_XNOR2 U105 ( .A(n95), .B(n93), .Z(sum[1]) );
  GTECH_AO22 U106 ( .A(n96), .B(cin), .C(a[0]), .D(b[0]), .Z(n93) );
  GTECH_NOT U107 ( .A(n94), .Z(n95) );
  GTECH_XNOR2 U108 ( .A(n97), .B(n98), .Z(sum[15]) );
  GTECH_OAI21 U109 ( .A(n99), .B(n100), .C(n101), .Z(n98) );
  GTECH_XOR2 U110 ( .A(n100), .B(n99), .Z(sum[14]) );
  GTECH_OA21 U111 ( .A(n102), .B(n103), .C(n104), .Z(n99) );
  GTECH_XOR2 U112 ( .A(n103), .B(n102), .Z(sum[13]) );
  GTECH_OA21 U113 ( .A(n105), .B(n106), .C(n107), .Z(n102) );
  GTECH_XOR2 U114 ( .A(n105), .B(n106), .Z(sum[12]) );
  GTECH_NOT U115 ( .A(cout), .Z(n105) );
  GTECH_XNOR2 U116 ( .A(n108), .B(n109), .Z(sum[11]) );
  GTECH_OAI21 U117 ( .A(n110), .B(n111), .C(n112), .Z(n108) );
  GTECH_XOR2 U118 ( .A(n110), .B(n111), .Z(sum[10]) );
  GTECH_OA21 U119 ( .A(n74), .B(n73), .C(n113), .Z(n110) );
  GTECH_OA21 U120 ( .A(n76), .B(n75), .C(n114), .Z(n74) );
  GTECH_NOT U121 ( .A(n115), .Z(n76) );
  GTECH_XNOR2 U122 ( .A(cin), .B(n116), .Z(sum[0]) );
  GTECH_AO21 U123 ( .A(n115), .B(n117), .C(n118), .Z(cout) );
  GTECH_AO21 U124 ( .A(n85), .B(n119), .C(n120), .Z(n115) );
  GTECH_NAND2 U125 ( .A(n121), .B(n122), .Z(n85) );
  GTECH_NAND4 U126 ( .A(n123), .B(n92), .C(cin), .D(n124), .Z(n122) );
  GTECH_AND3 U127 ( .A(n125), .B(n94), .C(n96), .Z(n124) );
  GTECH_AND4 U128 ( .A(n119), .B(n123), .C(n117), .D(n126), .Z(Pm) );
  GTECH_AND4 U129 ( .A(n92), .B(n96), .C(n125), .D(n94), .Z(n126) );
  GTECH_NOT U130 ( .A(n87), .Z(n125) );
  GTECH_NOT U131 ( .A(n116), .Z(n96) );
  GTECH_XNOR2 U132 ( .A(a[0]), .B(b[0]), .Z(n116) );
  GTECH_AO21 U133 ( .A(n127), .B(n117), .C(n118), .Z(Gm) );
  GTECH_OAI2N2 U134 ( .A(n128), .B(n97), .C(b[15]), .D(a[15]), .Z(n118) );
  GTECH_OA21 U135 ( .A(n129), .B(n100), .C(n101), .Z(n128) );
  GTECH_OA21 U136 ( .A(n107), .B(n103), .C(n104), .Z(n129) );
  GTECH_NOR4 U137 ( .A(n106), .B(n100), .C(n103), .D(n97), .Z(n117) );
  GTECH_XNOR2 U138 ( .A(a[15]), .B(b[15]), .Z(n97) );
  GTECH_OAI21 U139 ( .A(b[13]), .B(a[13]), .C(n104), .Z(n103) );
  GTECH_NAND2 U140 ( .A(b[13]), .B(a[13]), .Z(n104) );
  GTECH_OAI21 U141 ( .A(b[14]), .B(a[14]), .C(n101), .Z(n100) );
  GTECH_NAND2 U142 ( .A(b[14]), .B(a[14]), .Z(n101) );
  GTECH_OAI21 U143 ( .A(b[12]), .B(a[12]), .C(n107), .Z(n106) );
  GTECH_NAND2 U144 ( .A(b[12]), .B(a[12]), .Z(n107) );
  GTECH_AO21 U145 ( .A(n130), .B(n119), .C(n120), .Z(n127) );
  GTECH_OAI21 U146 ( .A(n131), .B(n109), .C(n132), .Z(n120) );
  GTECH_OA21 U147 ( .A(n133), .B(n111), .C(n112), .Z(n131) );
  GTECH_OA21 U148 ( .A(n73), .B(n114), .C(n113), .Z(n133) );
  GTECH_NAND2 U149 ( .A(a[9]), .B(b[9]), .Z(n113) );
  GTECH_NOR4 U150 ( .A(n75), .B(n109), .C(n111), .D(n73), .Z(n119) );
  GTECH_XNOR2 U151 ( .A(a[9]), .B(b[9]), .Z(n73) );
  GTECH_OAI21 U152 ( .A(a[10]), .B(b[10]), .C(n112), .Z(n111) );
  GTECH_NAND2 U153 ( .A(b[10]), .B(a[10]), .Z(n112) );
  GTECH_OAI21 U154 ( .A(a[11]), .B(b[11]), .C(n132), .Z(n109) );
  GTECH_NAND2 U155 ( .A(b[11]), .B(a[11]), .Z(n132) );
  GTECH_OAI21 U156 ( .A(b[8]), .B(a[8]), .C(n114), .Z(n75) );
  GTECH_NAND2 U157 ( .A(b[8]), .B(a[8]), .Z(n114) );
  GTECH_NOT U158 ( .A(n121), .Z(n130) );
  GTECH_AOI222 U159 ( .A(n123), .B(n134), .C(b[7]), .D(a[7]), .E(n77), .F(n135), .Z(n121) );
  GTECH_OAI21 U160 ( .A(n136), .B(n80), .C(n81), .Z(n135) );
  GTECH_NOT U161 ( .A(n82), .Z(n80) );
  GTECH_OA21 U162 ( .A(n137), .B(n138), .C(n139), .Z(n136) );
  GTECH_NAND3 U163 ( .A(a[4]), .B(n84), .C(b[4]), .Z(n139) );
  GTECH_NOT U164 ( .A(a[5]), .Z(n138) );
  GTECH_OAI2N2 U165 ( .A(n140), .B(n87), .C(b[3]), .D(a[3]), .Z(n134) );
  GTECH_XNOR2 U166 ( .A(a[3]), .B(b[3]), .Z(n87) );
  GTECH_OA21 U167 ( .A(n141), .B(n90), .C(n91), .Z(n140) );
  GTECH_NOT U168 ( .A(n92), .Z(n90) );
  GTECH_OA21 U169 ( .A(a[2]), .B(b[2]), .C(n91), .Z(n92) );
  GTECH_NAND2 U170 ( .A(b[2]), .B(a[2]), .Z(n91) );
  GTECH_OA21 U171 ( .A(n142), .B(n143), .C(n144), .Z(n141) );
  GTECH_NAND3 U172 ( .A(a[0]), .B(n94), .C(b[0]), .Z(n144) );
  GTECH_XNOR2 U173 ( .A(a[1]), .B(n142), .Z(n94) );
  GTECH_NOT U174 ( .A(a[1]), .Z(n143) );
  GTECH_NOT U175 ( .A(b[1]), .Z(n142) );
  GTECH_AND4 U176 ( .A(n82), .B(n86), .C(n84), .D(n77), .Z(n123) );
  GTECH_XOR2 U177 ( .A(a[7]), .B(b[7]), .Z(n77) );
  GTECH_XNOR2 U178 ( .A(a[5]), .B(n137), .Z(n84) );
  GTECH_NOT U179 ( .A(b[5]), .Z(n137) );
  GTECH_XOR2 U180 ( .A(a[4]), .B(b[4]), .Z(n86) );
  GTECH_OA21 U181 ( .A(a[6]), .B(b[6]), .C(n81), .Z(n82) );
  GTECH_NAND2 U182 ( .A(b[6]), .B(a[6]), .Z(n81) );
endmodule

