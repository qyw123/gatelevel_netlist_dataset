
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392;

  GTECH_MUX2 U135 ( .A(n274), .B(n275), .S(n276), .Z(sum[9]) );
  GTECH_XNOR2 U136 ( .A(n277), .B(n278), .Z(n275) );
  GTECH_XNOR2 U137 ( .A(n279), .B(n277), .Z(n274) );
  GTECH_AO21 U138 ( .A(n280), .B(n281), .C(n282), .Z(n277) );
  GTECH_NOT U139 ( .A(b[9]), .Z(n281) );
  GTECH_OR_NOT U140 ( .A(n283), .B(n284), .Z(sum[8]) );
  GTECH_OAI21 U141 ( .A(n278), .B(n285), .C(n286), .Z(n284) );
  GTECH_MUX2 U142 ( .A(n287), .B(n288), .S(n289), .Z(sum[7]) );
  GTECH_XNOR2 U143 ( .A(n290), .B(n291), .Z(n288) );
  GTECH_AND2 U144 ( .A(n292), .B(n293), .Z(n291) );
  GTECH_OAI21 U145 ( .A(b[6]), .B(a[6]), .C(n294), .Z(n293) );
  GTECH_XOR2 U146 ( .A(n290), .B(n295), .Z(n287) );
  GTECH_XOR2 U147 ( .A(a[7]), .B(b[7]), .Z(n290) );
  GTECH_OAI21 U148 ( .A(n296), .B(n292), .C(n297), .Z(sum[6]) );
  GTECH_MUX2 U149 ( .A(n298), .B(n299), .S(b[6]), .Z(n297) );
  GTECH_OR_NOT U150 ( .A(a[6]), .B(n296), .Z(n299) );
  GTECH_XOR2 U151 ( .A(a[6]), .B(n296), .Z(n298) );
  GTECH_NOT U152 ( .A(n300), .Z(n296) );
  GTECH_AO21 U153 ( .A(n301), .B(n302), .C(n294), .Z(n300) );
  GTECH_OA21 U154 ( .A(n303), .B(n304), .C(n305), .Z(n294) );
  GTECH_MUX2 U155 ( .A(n306), .B(n307), .S(n308), .Z(sum[5]) );
  GTECH_AND_NOT U156 ( .A(n305), .B(n304), .Z(n308) );
  GTECH_AO21 U157 ( .A(n309), .B(n289), .C(n310), .Z(n307) );
  GTECH_AO21 U158 ( .A(n311), .B(n301), .C(n303), .Z(n306) );
  GTECH_NOT U159 ( .A(n309), .Z(n303) );
  GTECH_XNOR2 U160 ( .A(n312), .B(n301), .Z(sum[4]) );
  GTECH_NOT U161 ( .A(n289), .Z(n301) );
  GTECH_MUX2 U162 ( .A(n313), .B(n314), .S(n315), .Z(sum[3]) );
  GTECH_XOR2 U163 ( .A(n316), .B(n317), .Z(n314) );
  GTECH_AO21 U164 ( .A(n318), .B(n319), .C(n320), .Z(n317) );
  GTECH_XOR2 U165 ( .A(n316), .B(n321), .Z(n313) );
  GTECH_XOR2 U166 ( .A(a[3]), .B(b[3]), .Z(n316) );
  GTECH_MUX2 U167 ( .A(n322), .B(n323), .S(cin), .Z(sum[2]) );
  GTECH_MUX2 U168 ( .A(n324), .B(n325), .S(n326), .Z(n323) );
  GTECH_MUX2 U169 ( .A(n324), .B(n325), .S(n319), .Z(n322) );
  GTECH_OA21 U170 ( .A(n327), .B(n328), .C(n329), .Z(n319) );
  GTECH_OR_NOT U171 ( .A(n320), .B(n318), .Z(n325) );
  GTECH_XOR2 U172 ( .A(a[2]), .B(b[2]), .Z(n324) );
  GTECH_MUX2 U173 ( .A(n330), .B(n331), .S(n332), .Z(sum[1]) );
  GTECH_AND_NOT U174 ( .A(n329), .B(n327), .Z(n332) );
  GTECH_AO21 U175 ( .A(n315), .B(n333), .C(n334), .Z(n331) );
  GTECH_AO21 U176 ( .A(n335), .B(cin), .C(n328), .Z(n330) );
  GTECH_NOT U177 ( .A(n333), .Z(n328) );
  GTECH_MUX2 U178 ( .A(n336), .B(n337), .S(n338), .Z(sum[15]) );
  GTECH_XNOR2 U179 ( .A(n339), .B(n340), .Z(n337) );
  GTECH_XNOR2 U180 ( .A(n339), .B(n341), .Z(n336) );
  GTECH_AND2 U181 ( .A(n342), .B(n343), .Z(n341) );
  GTECH_OAI21 U182 ( .A(b[14]), .B(a[14]), .C(n344), .Z(n343) );
  GTECH_XOR2 U183 ( .A(a[15]), .B(b[15]), .Z(n339) );
  GTECH_OAI21 U184 ( .A(n345), .B(n342), .C(n346), .Z(sum[14]) );
  GTECH_MUX2 U185 ( .A(n347), .B(n348), .S(b[14]), .Z(n346) );
  GTECH_OR_NOT U186 ( .A(a[14]), .B(n345), .Z(n348) );
  GTECH_XOR2 U187 ( .A(a[14]), .B(n345), .Z(n347) );
  GTECH_NOT U188 ( .A(n349), .Z(n345) );
  GTECH_AO21 U189 ( .A(n338), .B(n350), .C(n344), .Z(n349) );
  GTECH_OAI21 U190 ( .A(n351), .B(n352), .C(n353), .Z(n344) );
  GTECH_MUX2 U191 ( .A(n354), .B(n355), .S(n356), .Z(sum[13]) );
  GTECH_OA21 U192 ( .A(n357), .B(n358), .C(n352), .Z(n356) );
  GTECH_XOR2 U193 ( .A(b[13]), .B(a[13]), .Z(n355) );
  GTECH_OR_NOT U194 ( .A(n351), .B(n353), .Z(n354) );
  GTECH_NAND2 U195 ( .A(n359), .B(n360), .Z(sum[12]) );
  GTECH_AO21 U196 ( .A(n352), .B(n361), .C(n357), .Z(n359) );
  GTECH_MUX2 U197 ( .A(n362), .B(n363), .S(n276), .Z(sum[11]) );
  GTECH_XOR2 U198 ( .A(n364), .B(n365), .Z(n363) );
  GTECH_AO21 U199 ( .A(n366), .B(n367), .C(n368), .Z(n365) );
  GTECH_XOR2 U200 ( .A(n364), .B(n369), .Z(n362) );
  GTECH_XOR2 U201 ( .A(a[11]), .B(b[11]), .Z(n364) );
  GTECH_MUX2 U202 ( .A(n370), .B(n371), .S(n372), .Z(sum[10]) );
  GTECH_OA21 U203 ( .A(n367), .B(n286), .C(n373), .Z(n372) );
  GTECH_OA21 U204 ( .A(n282), .B(n278), .C(n374), .Z(n367) );
  GTECH_OR_NOT U205 ( .A(n368), .B(n366), .Z(n371) );
  GTECH_XOR2 U206 ( .A(b[10]), .B(a[10]), .Z(n370) );
  GTECH_XNOR2 U207 ( .A(cin), .B(n375), .Z(sum[0]) );
  GTECH_OAI21 U208 ( .A(n357), .B(n376), .C(n360), .Z(cout) );
  GTECH_NAND3 U209 ( .A(n352), .B(n361), .C(n357), .Z(n360) );
  GTECH_NAND2 U210 ( .A(a[12]), .B(b[12]), .Z(n352) );
  GTECH_OA21 U211 ( .A(n340), .B(n377), .C(n378), .Z(n376) );
  GTECH_OAI21 U212 ( .A(a[15]), .B(n379), .C(b[15]), .Z(n378) );
  GTECH_NOT U213 ( .A(a[15]), .Z(n377) );
  GTECH_NOT U214 ( .A(n379), .Z(n340) );
  GTECH_NAND2 U215 ( .A(n380), .B(n342), .Z(n379) );
  GTECH_NAND2 U216 ( .A(b[14]), .B(a[14]), .Z(n342) );
  GTECH_OAI21 U217 ( .A(a[14]), .B(b[14]), .C(n350), .Z(n380) );
  GTECH_OAI21 U218 ( .A(n358), .B(n351), .C(n353), .Z(n350) );
  GTECH_NAND2 U219 ( .A(b[13]), .B(a[13]), .Z(n353) );
  GTECH_NOT U220 ( .A(n381), .Z(n351) );
  GTECH_OR2 U221 ( .A(a[13]), .B(b[13]), .Z(n381) );
  GTECH_NOT U222 ( .A(n361), .Z(n358) );
  GTECH_OR2 U223 ( .A(b[12]), .B(a[12]), .Z(n361) );
  GTECH_NOT U224 ( .A(n338), .Z(n357) );
  GTECH_AO21 U225 ( .A(n382), .B(n286), .C(n283), .Z(n338) );
  GTECH_NOR3 U226 ( .A(n278), .B(n285), .C(n286), .Z(n283) );
  GTECH_NOT U227 ( .A(n279), .Z(n285) );
  GTECH_AND2 U228 ( .A(b[8]), .B(a[8]), .Z(n278) );
  GTECH_NOT U229 ( .A(n276), .Z(n286) );
  GTECH_MUX2 U230 ( .A(n383), .B(n312), .S(n289), .Z(n276) );
  GTECH_MUX2 U231 ( .A(n384), .B(n375), .S(n315), .Z(n289) );
  GTECH_NOT U232 ( .A(cin), .Z(n315) );
  GTECH_OR_NOT U233 ( .A(n334), .B(n333), .Z(n375) );
  GTECH_NAND2 U234 ( .A(b[0]), .B(a[0]), .Z(n333) );
  GTECH_NOT U235 ( .A(n335), .Z(n334) );
  GTECH_NOT U236 ( .A(n385), .Z(n384) );
  GTECH_AO21 U237 ( .A(n321), .B(a[3]), .C(n386), .Z(n385) );
  GTECH_OA21 U238 ( .A(a[3]), .B(n321), .C(b[3]), .Z(n386) );
  GTECH_AO21 U239 ( .A(n318), .B(n326), .C(n320), .Z(n321) );
  GTECH_AND2 U240 ( .A(b[2]), .B(a[2]), .Z(n320) );
  GTECH_OA21 U241 ( .A(n327), .B(n335), .C(n329), .Z(n326) );
  GTECH_OR2 U242 ( .A(a[1]), .B(b[1]), .Z(n329) );
  GTECH_OR2 U243 ( .A(a[0]), .B(b[0]), .Z(n335) );
  GTECH_AND2 U244 ( .A(b[1]), .B(a[1]), .Z(n327) );
  GTECH_OR2 U245 ( .A(b[2]), .B(a[2]), .Z(n318) );
  GTECH_OR_NOT U246 ( .A(n310), .B(n309), .Z(n312) );
  GTECH_NAND2 U247 ( .A(b[4]), .B(a[4]), .Z(n309) );
  GTECH_NOT U248 ( .A(n311), .Z(n310) );
  GTECH_OA21 U249 ( .A(n387), .B(n388), .C(n389), .Z(n383) );
  GTECH_OAI21 U250 ( .A(a[7]), .B(n295), .C(b[7]), .Z(n389) );
  GTECH_NOT U251 ( .A(n387), .Z(n295) );
  GTECH_NOT U252 ( .A(a[7]), .Z(n388) );
  GTECH_AND2 U253 ( .A(n390), .B(n292), .Z(n387) );
  GTECH_NAND2 U254 ( .A(b[6]), .B(a[6]), .Z(n292) );
  GTECH_OAI21 U255 ( .A(a[6]), .B(b[6]), .C(n302), .Z(n390) );
  GTECH_OA21 U256 ( .A(n304), .B(n311), .C(n305), .Z(n302) );
  GTECH_OR2 U257 ( .A(b[5]), .B(a[5]), .Z(n305) );
  GTECH_OR2 U258 ( .A(a[4]), .B(b[4]), .Z(n311) );
  GTECH_AND2 U259 ( .A(a[5]), .B(b[5]), .Z(n304) );
  GTECH_AO21 U260 ( .A(n369), .B(a[11]), .C(n391), .Z(n382) );
  GTECH_OA21 U261 ( .A(a[11]), .B(n369), .C(b[11]), .Z(n391) );
  GTECH_AO21 U262 ( .A(n366), .B(n373), .C(n368), .Z(n369) );
  GTECH_AND_NOT U263 ( .A(b[10]), .B(n392), .Z(n368) );
  GTECH_NOT U264 ( .A(a[10]), .Z(n392) );
  GTECH_OA21 U265 ( .A(n282), .B(n279), .C(n374), .Z(n373) );
  GTECH_OR_NOT U266 ( .A(b[9]), .B(n280), .Z(n374) );
  GTECH_NOT U267 ( .A(a[9]), .Z(n280) );
  GTECH_OR2 U268 ( .A(a[8]), .B(b[8]), .Z(n279) );
  GTECH_AND2 U269 ( .A(a[9]), .B(b[9]), .Z(n282) );
  GTECH_OR2 U270 ( .A(b[10]), .B(a[10]), .Z(n366) );
endmodule

