
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135;

  GTECH_ADD_AB U87 ( .A(n68), .B(n69), .S(sum[9]) );
  GTECH_ADD_AB U88 ( .A(n70), .B(n71), .S(sum[8]) );
  GTECH_ADD_AB U89 ( .A(n72), .B(n73), .S(sum[7]) );
  GTECH_OA21 U90 ( .A(n74), .B(n75), .C(n76), .Z(n73) );
  GTECH_ADD_AB U91 ( .A(n74), .B(n75), .S(sum[6]) );
  GTECH_OA21 U92 ( .A(n77), .B(n78), .C(n79), .Z(n74) );
  GTECH_ADD_AB U93 ( .A(n77), .B(n78), .S(sum[5]) );
  GTECH_OA21 U94 ( .A(n80), .B(n81), .C(n82), .Z(n77) );
  GTECH_NOT U95 ( .A(n83), .Z(n80) );
  GTECH_XNOR2 U96 ( .A(n83), .B(n81), .Z(sum[4]) );
  GTECH_ADD_AB U97 ( .A(n84), .B(n85), .S(sum[3]) );
  GTECH_OA21 U98 ( .A(n86), .B(n87), .C(n88), .Z(n84) );
  GTECH_ADD_AB U99 ( .A(n86), .B(n87), .S(sum[2]) );
  GTECH_OA21 U100 ( .A(n89), .B(n90), .C(n91), .Z(n86) );
  GTECH_ADD_AB U101 ( .A(n89), .B(n90), .S(sum[1]) );
  GTECH_AND2 U102 ( .A(n92), .B(n93), .Z(n89) );
  GTECH_ADD_AB U103 ( .A(n94), .B(n95), .S(sum[15]) );
  GTECH_OA21 U104 ( .A(n96), .B(n97), .C(n98), .Z(n94) );
  GTECH_ADD_AB U105 ( .A(n96), .B(n97), .S(sum[14]) );
  GTECH_OA21 U106 ( .A(n99), .B(n100), .C(n101), .Z(n96) );
  GTECH_ADD_AB U107 ( .A(n99), .B(n100), .S(sum[13]) );
  GTECH_OA21 U108 ( .A(n102), .B(n103), .C(n104), .Z(n99) );
  GTECH_NOT U109 ( .A(cout), .Z(n102) );
  GTECH_XNOR2 U110 ( .A(n103), .B(cout), .Z(sum[12]) );
  GTECH_ADD_AB U111 ( .A(n105), .B(n106), .S(sum[11]) );
  GTECH_OA21 U112 ( .A(n107), .B(n108), .C(n109), .Z(n106) );
  GTECH_ADD_AB U113 ( .A(n107), .B(n108), .S(sum[10]) );
  GTECH_OA21 U114 ( .A(n68), .B(n69), .C(n110), .Z(n107) );
  GTECH_OA21 U115 ( .A(n70), .B(n71), .C(n111), .Z(n68) );
  GTECH_ADD_AB U116 ( .A(cin), .B(n112), .S(sum[0]) );
  GTECH_OAI21 U117 ( .A(n70), .B(n113), .C(n114), .Z(cout) );
  GTECH_AOI21 U118 ( .A(n83), .B(n115), .C(n116), .Z(n70) );
  GTECH_OR_NOT U119 ( .A(n117), .B(n118), .Z(n83) );
  GTECH_OR5 U120 ( .A(n90), .B(n85), .C(n87), .D(n92), .E(n119), .Z(n118) );
  GTECH_OR_NOT U121 ( .A(n120), .B(cin), .Z(n92) );
  GTECH_NOR4 U122 ( .A(n121), .B(n113), .C(n120), .D(n122), .Z(Pm) );
  GTECH_NOT U123 ( .A(n112), .Z(n120) );
  GTECH_OA21 U124 ( .A(b[0]), .B(a[0]), .C(n93), .Z(n112) );
  GTECH_OR4 U125 ( .A(n119), .B(n87), .C(n90), .D(n85), .Z(n121) );
  GTECH_OAI21 U126 ( .A(n123), .B(n113), .C(n114), .Z(Gm) );
  GTECH_AOI2N2 U127 ( .A(b[15]), .B(a[15]), .C(n124), .D(n95), .Z(n114) );
  GTECH_OA21 U128 ( .A(n125), .B(n97), .C(n98), .Z(n124) );
  GTECH_OA21 U129 ( .A(n104), .B(n100), .C(n101), .Z(n125) );
  GTECH_OR4 U130 ( .A(n103), .B(n97), .C(n100), .D(n95), .Z(n113) );
  GTECH_XNOR2 U131 ( .A(b[15]), .B(a[15]), .Z(n95) );
  GTECH_OAI21 U132 ( .A(b[13]), .B(a[13]), .C(n101), .Z(n100) );
  GTECH_NAND2 U133 ( .A(b[13]), .B(a[13]), .Z(n101) );
  GTECH_OAI21 U134 ( .A(b[14]), .B(a[14]), .C(n98), .Z(n97) );
  GTECH_NAND2 U135 ( .A(b[14]), .B(a[14]), .Z(n98) );
  GTECH_OAI21 U136 ( .A(b[12]), .B(a[12]), .C(n104), .Z(n103) );
  GTECH_NAND2 U137 ( .A(a[12]), .B(b[12]), .Z(n104) );
  GTECH_AOI21 U138 ( .A(n117), .B(n115), .C(n116), .Z(n123) );
  GTECH_OAI21 U139 ( .A(n126), .B(n105), .C(n127), .Z(n116) );
  GTECH_OA21 U140 ( .A(n128), .B(n108), .C(n109), .Z(n126) );
  GTECH_OA21 U141 ( .A(n111), .B(n69), .C(n110), .Z(n128) );
  GTECH_NOT U142 ( .A(n122), .Z(n115) );
  GTECH_OR4 U143 ( .A(n71), .B(n105), .C(n108), .D(n69), .Z(n122) );
  GTECH_OAI21 U144 ( .A(b[9]), .B(a[9]), .C(n110), .Z(n69) );
  GTECH_NAND2 U145 ( .A(b[9]), .B(a[9]), .Z(n110) );
  GTECH_OAI21 U146 ( .A(b[10]), .B(a[10]), .C(n109), .Z(n108) );
  GTECH_NAND2 U147 ( .A(b[10]), .B(a[10]), .Z(n109) );
  GTECH_OAI21 U148 ( .A(b[11]), .B(a[11]), .C(n127), .Z(n105) );
  GTECH_NAND2 U149 ( .A(a[11]), .B(b[11]), .Z(n127) );
  GTECH_OAI21 U150 ( .A(b[8]), .B(a[8]), .C(n111), .Z(n71) );
  GTECH_NAND2 U151 ( .A(a[8]), .B(b[8]), .Z(n111) );
  GTECH_OAI21 U152 ( .A(n129), .B(n119), .C(n130), .Z(n117) );
  GTECH_OA21 U153 ( .A(n131), .B(n72), .C(n132), .Z(n130) );
  GTECH_OA21 U154 ( .A(n133), .B(n75), .C(n76), .Z(n131) );
  GTECH_OA21 U155 ( .A(n78), .B(n82), .C(n79), .Z(n133) );
  GTECH_OR4 U156 ( .A(n81), .B(n72), .C(n75), .D(n78), .Z(n119) );
  GTECH_OAI21 U157 ( .A(b[5]), .B(a[5]), .C(n79), .Z(n78) );
  GTECH_NAND2 U158 ( .A(b[5]), .B(a[5]), .Z(n79) );
  GTECH_OAI21 U159 ( .A(b[6]), .B(a[6]), .C(n76), .Z(n75) );
  GTECH_NAND2 U160 ( .A(b[6]), .B(a[6]), .Z(n76) );
  GTECH_OAI21 U161 ( .A(b[7]), .B(a[7]), .C(n132), .Z(n72) );
  GTECH_NAND2 U162 ( .A(a[7]), .B(b[7]), .Z(n132) );
  GTECH_OAI21 U163 ( .A(b[4]), .B(a[4]), .C(n82), .Z(n81) );
  GTECH_NAND2 U164 ( .A(a[4]), .B(b[4]), .Z(n82) );
  GTECH_AOI2N2 U165 ( .A(b[3]), .B(a[3]), .C(n134), .D(n85), .Z(n129) );
  GTECH_XNOR2 U166 ( .A(b[3]), .B(a[3]), .Z(n85) );
  GTECH_OA21 U167 ( .A(n135), .B(n87), .C(n88), .Z(n134) );
  GTECH_OAI21 U168 ( .A(b[2]), .B(a[2]), .C(n88), .Z(n87) );
  GTECH_NAND2 U169 ( .A(b[2]), .B(a[2]), .Z(n88) );
  GTECH_OA21 U170 ( .A(n90), .B(n93), .C(n91), .Z(n135) );
  GTECH_NAND2 U171 ( .A(b[0]), .B(a[0]), .Z(n93) );
  GTECH_OAI21 U172 ( .A(b[1]), .B(a[1]), .C(n91), .Z(n90) );
  GTECH_NAND2 U173 ( .A(b[1]), .B(a[1]), .Z(n91) );
endmodule

