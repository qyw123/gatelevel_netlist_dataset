
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_OAI21 U75 ( .A(n83), .B(n84), .C(n85), .Z(N155) );
  GTECH_OA22 U76 ( .A(n86), .B(n87), .C(n88), .D(n89), .Z(n85) );
  GTECH_NOT U77 ( .A(n90), .Z(n87) );
  GTECH_XOR2 U78 ( .A(n91), .B(n92), .Z(N154) );
  GTECH_NOT U79 ( .A(n83), .Z(n92) );
  GTECH_XOR2 U80 ( .A(n90), .B(n86), .Z(n83) );
  GTECH_AOI2N2 U81 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n86) );
  GTECH_OR_NOT U82 ( .A(n97), .B(n95), .Z(n94) );
  GTECH_XOR2 U83 ( .A(n89), .B(n88), .Z(n90) );
  GTECH_AND2 U84 ( .A(n98), .B(n99), .Z(n88) );
  GTECH_OR_NOT U85 ( .A(n100), .B(n101), .Z(n99) );
  GTECH_OAI21 U86 ( .A(n102), .B(n101), .C(n103), .Z(n98) );
  GTECH_OR_NOT U87 ( .A(n104), .B(I_b[7]), .Z(n89) );
  GTECH_NOT U88 ( .A(n84), .Z(n91) );
  GTECH_OR_NOT U89 ( .A(n105), .B(n106), .Z(n84) );
  GTECH_XOR2 U90 ( .A(n107), .B(n106), .Z(N153) );
  GTECH_NOT U91 ( .A(n108), .Z(n106) );
  GTECH_XOR3 U92 ( .A(n97), .B(n95), .C(n93), .Z(n108) );
  GTECH_XOR3 U93 ( .A(n102), .B(n103), .C(n101), .Z(n93) );
  GTECH_OAI21 U94 ( .A(n109), .B(n110), .C(n111), .Z(n101) );
  GTECH_OAI21 U95 ( .A(n112), .B(n113), .C(n114), .Z(n111) );
  GTECH_NOT U96 ( .A(n113), .Z(n109) );
  GTECH_NOT U97 ( .A(n115), .Z(n103) );
  GTECH_OR_NOT U98 ( .A(n116), .B(I_b[7]), .Z(n115) );
  GTECH_NOT U99 ( .A(n100), .Z(n102) );
  GTECH_OR_NOT U100 ( .A(n117), .B(I_a[7]), .Z(n100) );
  GTECH_NOT U101 ( .A(I_b[6]), .Z(n117) );
  GTECH_ADD_ABC U102 ( .A(n118), .B(n119), .C(n120), .COUT(n95) );
  GTECH_NOT U103 ( .A(n121), .Z(n120) );
  GTECH_XOR2 U104 ( .A(n122), .B(n123), .Z(n119) );
  GTECH_AND2 U105 ( .A(I_a[7]), .B(I_b[5]), .Z(n123) );
  GTECH_NOT U106 ( .A(n96), .Z(n97) );
  GTECH_OR_NOT U107 ( .A(n122), .B(I_a[7]), .Z(n96) );
  GTECH_NOT U108 ( .A(n105), .Z(n107) );
  GTECH_OR_NOT U109 ( .A(n124), .B(n125), .Z(n105) );
  GTECH_XOR2 U110 ( .A(n124), .B(n126), .Z(N152) );
  GTECH_NOT U111 ( .A(n125), .Z(n126) );
  GTECH_XOR4 U112 ( .A(n127), .B(n122), .C(n118), .D(n121), .Z(n125) );
  GTECH_XOR3 U113 ( .A(n112), .B(n114), .C(n113), .Z(n121) );
  GTECH_OAI21 U114 ( .A(n128), .B(n129), .C(n130), .Z(n113) );
  GTECH_OAI21 U115 ( .A(n131), .B(n132), .C(n133), .Z(n130) );
  GTECH_NOT U116 ( .A(n132), .Z(n128) );
  GTECH_NOT U117 ( .A(n134), .Z(n114) );
  GTECH_OR_NOT U118 ( .A(n135), .B(I_b[7]), .Z(n134) );
  GTECH_NOT U119 ( .A(n110), .Z(n112) );
  GTECH_OR_NOT U120 ( .A(n116), .B(I_b[6]), .Z(n110) );
  GTECH_NOT U121 ( .A(I_a[6]), .Z(n116) );
  GTECH_ADD_ABC U122 ( .A(n136), .B(n137), .C(n138), .COUT(n118) );
  GTECH_NOT U123 ( .A(n139), .Z(n138) );
  GTECH_XOR3 U124 ( .A(n140), .B(n141), .C(n142), .Z(n137) );
  GTECH_OA21 U125 ( .A(n142), .B(n143), .C(n144), .Z(n122) );
  GTECH_OAI21 U126 ( .A(n140), .B(n145), .C(n141), .Z(n144) );
  GTECH_NOT U127 ( .A(n143), .Z(n140) );
  GTECH_NOT U128 ( .A(n145), .Z(n142) );
  GTECH_AND2 U129 ( .A(I_b[5]), .B(I_a[7]), .Z(n127) );
  GTECH_ADD_ABC U130 ( .A(n146), .B(n147), .C(n148), .COUT(n124) );
  GTECH_NOT U131 ( .A(n149), .Z(n148) );
  GTECH_OA22 U132 ( .A(n150), .B(n104), .C(n151), .D(n152), .Z(n147) );
  GTECH_OA21 U133 ( .A(n153), .B(n154), .C(n155), .Z(n146) );
  GTECH_XOR3 U134 ( .A(n156), .B(n149), .C(n157), .Z(N151) );
  GTECH_OA21 U135 ( .A(n153), .B(n154), .C(n155), .Z(n157) );
  GTECH_OAI21 U136 ( .A(n158), .B(n159), .C(n160), .Z(n155) );
  GTECH_XOR2 U137 ( .A(n161), .B(n136), .Z(n149) );
  GTECH_ADD_ABC U138 ( .A(n162), .B(n163), .C(n164), .COUT(n136) );
  GTECH_NOT U139 ( .A(n165), .Z(n164) );
  GTECH_XOR3 U140 ( .A(n166), .B(n167), .C(n168), .Z(n163) );
  GTECH_XOR4 U141 ( .A(n141), .B(n145), .C(n143), .D(n139), .Z(n161) );
  GTECH_XOR3 U142 ( .A(n131), .B(n133), .C(n132), .Z(n139) );
  GTECH_OAI21 U143 ( .A(n169), .B(n170), .C(n171), .Z(n132) );
  GTECH_OAI21 U144 ( .A(n172), .B(n173), .C(n174), .Z(n171) );
  GTECH_NOT U145 ( .A(n173), .Z(n169) );
  GTECH_NOT U146 ( .A(n175), .Z(n133) );
  GTECH_OR_NOT U147 ( .A(n176), .B(I_b[7]), .Z(n175) );
  GTECH_NOT U148 ( .A(n129), .Z(n131) );
  GTECH_OR_NOT U149 ( .A(n135), .B(I_b[6]), .Z(n129) );
  GTECH_NOT U150 ( .A(I_a[5]), .Z(n135) );
  GTECH_OR_NOT U151 ( .A(n177), .B(I_a[7]), .Z(n143) );
  GTECH_OAI21 U152 ( .A(n168), .B(n178), .C(n179), .Z(n145) );
  GTECH_OAI21 U153 ( .A(n166), .B(n180), .C(n167), .Z(n179) );
  GTECH_NOT U154 ( .A(n178), .Z(n166) );
  GTECH_NOT U155 ( .A(n180), .Z(n168) );
  GTECH_NOT U156 ( .A(n181), .Z(n141) );
  GTECH_OR_NOT U157 ( .A(n182), .B(I_a[6]), .Z(n181) );
  GTECH_OA22 U158 ( .A(n150), .B(n104), .C(n151), .D(n152), .Z(n156) );
  GTECH_NOT U159 ( .A(n183), .Z(n152) );
  GTECH_NOT U160 ( .A(I_a[7]), .Z(n104) );
  GTECH_XOR3 U161 ( .A(n153), .B(n158), .C(n184), .Z(N150) );
  GTECH_NOT U162 ( .A(n160), .Z(n184) );
  GTECH_XOR2 U163 ( .A(n185), .B(n162), .Z(n160) );
  GTECH_ADD_ABC U164 ( .A(n186), .B(n187), .C(n188), .COUT(n162) );
  GTECH_NOT U165 ( .A(n189), .Z(n188) );
  GTECH_XOR3 U166 ( .A(n190), .B(n191), .C(n192), .Z(n187) );
  GTECH_XOR4 U167 ( .A(n167), .B(n180), .C(n178), .D(n165), .Z(n185) );
  GTECH_XOR3 U168 ( .A(n172), .B(n174), .C(n173), .Z(n165) );
  GTECH_OAI21 U169 ( .A(n193), .B(n194), .C(n195), .Z(n173) );
  GTECH_OAI21 U170 ( .A(n196), .B(n197), .C(n198), .Z(n195) );
  GTECH_NOT U171 ( .A(n197), .Z(n193) );
  GTECH_NOT U172 ( .A(n199), .Z(n174) );
  GTECH_OR_NOT U173 ( .A(n200), .B(I_b[7]), .Z(n199) );
  GTECH_NOT U174 ( .A(n170), .Z(n172) );
  GTECH_OR_NOT U175 ( .A(n176), .B(I_b[6]), .Z(n170) );
  GTECH_OR_NOT U176 ( .A(n177), .B(I_a[6]), .Z(n178) );
  GTECH_OAI21 U177 ( .A(n192), .B(n201), .C(n202), .Z(n180) );
  GTECH_OAI21 U178 ( .A(n190), .B(n203), .C(n191), .Z(n202) );
  GTECH_NOT U179 ( .A(n201), .Z(n190) );
  GTECH_NOT U180 ( .A(n203), .Z(n192) );
  GTECH_NOT U181 ( .A(n204), .Z(n167) );
  GTECH_OR_NOT U182 ( .A(n182), .B(I_a[5]), .Z(n204) );
  GTECH_NOT U183 ( .A(I_b[5]), .Z(n182) );
  GTECH_NOT U184 ( .A(n154), .Z(n158) );
  GTECH_XOR2 U185 ( .A(n183), .B(n151), .Z(n154) );
  GTECH_AOI2N2 U186 ( .A(n205), .B(n206), .C(n207), .D(n208), .Z(n151) );
  GTECH_OR_NOT U187 ( .A(n209), .B(n207), .Z(n206) );
  GTECH_XOR2 U188 ( .A(n210), .B(n150), .Z(n183) );
  GTECH_AND2 U189 ( .A(n211), .B(n212), .Z(n150) );
  GTECH_OR_NOT U190 ( .A(n213), .B(n214), .Z(n212) );
  GTECH_OAI21 U191 ( .A(n215), .B(n214), .C(n216), .Z(n211) );
  GTECH_OR_NOT U192 ( .A(n217), .B(I_a[7]), .Z(n210) );
  GTECH_NOT U193 ( .A(n159), .Z(n153) );
  GTECH_OAI2N2 U194 ( .A(n218), .B(n219), .C(n220), .D(n221), .Z(n159) );
  GTECH_OR_NOT U195 ( .A(n222), .B(n218), .Z(n221) );
  GTECH_XOR3 U196 ( .A(n218), .B(n222), .C(n223), .Z(N149) );
  GTECH_NOT U197 ( .A(n220), .Z(n223) );
  GTECH_XOR2 U198 ( .A(n224), .B(n186), .Z(n220) );
  GTECH_ADD_ABC U199 ( .A(n225), .B(n226), .C(n227), .COUT(n186) );
  GTECH_XOR3 U200 ( .A(n228), .B(n229), .C(n230), .Z(n226) );
  GTECH_OA21 U201 ( .A(n231), .B(n232), .C(n233), .Z(n225) );
  GTECH_XOR4 U202 ( .A(n191), .B(n203), .C(n201), .D(n189), .Z(n224) );
  GTECH_XOR3 U203 ( .A(n196), .B(n198), .C(n197), .Z(n189) );
  GTECH_OAI21 U204 ( .A(n234), .B(n235), .C(n236), .Z(n197) );
  GTECH_NOT U205 ( .A(n237), .Z(n198) );
  GTECH_OR_NOT U206 ( .A(n238), .B(I_b[7]), .Z(n237) );
  GTECH_NOT U207 ( .A(n194), .Z(n196) );
  GTECH_OR_NOT U208 ( .A(n200), .B(I_b[6]), .Z(n194) );
  GTECH_OR_NOT U209 ( .A(n177), .B(I_a[5]), .Z(n201) );
  GTECH_NOT U210 ( .A(I_b[4]), .Z(n177) );
  GTECH_OAI21 U211 ( .A(n230), .B(n239), .C(n240), .Z(n203) );
  GTECH_OAI21 U212 ( .A(n228), .B(n241), .C(n229), .Z(n240) );
  GTECH_NOT U213 ( .A(n239), .Z(n228) );
  GTECH_NOT U214 ( .A(n241), .Z(n230) );
  GTECH_NOT U215 ( .A(n242), .Z(n191) );
  GTECH_OR_NOT U216 ( .A(n176), .B(I_b[5]), .Z(n242) );
  GTECH_NOT U217 ( .A(n219), .Z(n222) );
  GTECH_XOR3 U218 ( .A(n209), .B(n207), .C(n205), .Z(n219) );
  GTECH_XOR3 U219 ( .A(n215), .B(n216), .C(n214), .Z(n205) );
  GTECH_OAI21 U220 ( .A(n243), .B(n244), .C(n245), .Z(n214) );
  GTECH_OAI21 U221 ( .A(n246), .B(n247), .C(n248), .Z(n245) );
  GTECH_NOT U222 ( .A(n247), .Z(n243) );
  GTECH_NOT U223 ( .A(n249), .Z(n216) );
  GTECH_OR_NOT U224 ( .A(n217), .B(I_a[6]), .Z(n249) );
  GTECH_NOT U225 ( .A(n213), .Z(n215) );
  GTECH_OR_NOT U226 ( .A(n250), .B(I_a[7]), .Z(n213) );
  GTECH_ADD_ABC U227 ( .A(n251), .B(n252), .C(n253), .COUT(n207) );
  GTECH_XOR2 U228 ( .A(n254), .B(n255), .Z(n252) );
  GTECH_AND2 U229 ( .A(I_a[7]), .B(I_b[1]), .Z(n255) );
  GTECH_NOT U230 ( .A(n208), .Z(n209) );
  GTECH_OR_NOT U231 ( .A(n254), .B(I_a[7]), .Z(n208) );
  GTECH_ADD_ABC U232 ( .A(n256), .B(n257), .C(n258), .COUT(n218) );
  GTECH_XOR3 U233 ( .A(n251), .B(n259), .C(n253), .Z(n257) );
  GTECH_NOT U234 ( .A(n260), .Z(n253) );
  GTECH_XOR2 U235 ( .A(n256), .B(n261), .Z(N148) );
  GTECH_XOR4 U236 ( .A(n259), .B(n260), .C(n258), .D(n251), .Z(n261) );
  GTECH_ADD_ABC U237 ( .A(n262), .B(n263), .C(n264), .COUT(n251) );
  GTECH_XOR3 U238 ( .A(n265), .B(n266), .C(n267), .Z(n263) );
  GTECH_XOR2 U239 ( .A(n268), .B(n269), .Z(n258) );
  GTECH_OA21 U240 ( .A(n231), .B(n232), .C(n233), .Z(n269) );
  GTECH_OAI21 U241 ( .A(n270), .B(n271), .C(n272), .Z(n233) );
  GTECH_NOT U242 ( .A(n231), .Z(n271) );
  GTECH_XOR4 U243 ( .A(n229), .B(n241), .C(n239), .D(n227), .Z(n268) );
  GTECH_XOR3 U244 ( .A(n273), .B(n274), .C(n236), .Z(n227) );
  GTECH_NAND3 U245 ( .A(I_b[6]), .B(I_a[1]), .C(n275), .Z(n236) );
  GTECH_NOT U246 ( .A(n235), .Z(n274) );
  GTECH_OR_NOT U247 ( .A(n276), .B(I_b[7]), .Z(n235) );
  GTECH_NOT U248 ( .A(n234), .Z(n273) );
  GTECH_OR_NOT U249 ( .A(n238), .B(I_b[6]), .Z(n234) );
  GTECH_OR_NOT U250 ( .A(n176), .B(I_b[4]), .Z(n239) );
  GTECH_OAI21 U251 ( .A(n277), .B(n278), .C(n279), .Z(n241) );
  GTECH_OAI21 U252 ( .A(n280), .B(n281), .C(n282), .Z(n279) );
  GTECH_NOT U253 ( .A(n281), .Z(n277) );
  GTECH_NOT U254 ( .A(n283), .Z(n229) );
  GTECH_OR_NOT U255 ( .A(n200), .B(I_b[5]), .Z(n283) );
  GTECH_XOR3 U256 ( .A(n246), .B(n248), .C(n247), .Z(n260) );
  GTECH_OAI21 U257 ( .A(n284), .B(n285), .C(n286), .Z(n247) );
  GTECH_OAI21 U258 ( .A(n287), .B(n288), .C(n289), .Z(n286) );
  GTECH_NOT U259 ( .A(n288), .Z(n284) );
  GTECH_NOT U260 ( .A(n290), .Z(n248) );
  GTECH_OR_NOT U261 ( .A(n217), .B(I_a[5]), .Z(n290) );
  GTECH_NOT U262 ( .A(I_b[3]), .Z(n217) );
  GTECH_NOT U263 ( .A(n244), .Z(n246) );
  GTECH_OR_NOT U264 ( .A(n250), .B(I_a[6]), .Z(n244) );
  GTECH_XOR2 U265 ( .A(n291), .B(n254), .Z(n259) );
  GTECH_OA21 U266 ( .A(n267), .B(n292), .C(n293), .Z(n254) );
  GTECH_OAI21 U267 ( .A(n265), .B(n294), .C(n266), .Z(n293) );
  GTECH_NOT U268 ( .A(n294), .Z(n267) );
  GTECH_AND2 U269 ( .A(I_b[1]), .B(I_a[7]), .Z(n291) );
  GTECH_ADD_ABC U270 ( .A(n295), .B(n296), .C(n297), .COUT(n256) );
  GTECH_NOT U271 ( .A(n298), .Z(n297) );
  GTECH_XOR3 U272 ( .A(n262), .B(n299), .C(n264), .Z(n296) );
  GTECH_NOT U273 ( .A(n300), .Z(n264) );
  GTECH_NOT U274 ( .A(n301), .Z(n299) );
  GTECH_XOR2 U275 ( .A(n302), .B(n295), .Z(N147) );
  GTECH_ADD_ABC U276 ( .A(n303), .B(n304), .C(n305), .COUT(n295) );
  GTECH_XOR3 U277 ( .A(n306), .B(n307), .C(n308), .Z(n304) );
  GTECH_OA21 U278 ( .A(n309), .B(n310), .C(n311), .Z(n303) );
  GTECH_XOR4 U279 ( .A(n300), .B(n262), .C(n301), .D(n298), .Z(n302) );
  GTECH_XOR3 U280 ( .A(n272), .B(n232), .C(n231), .Z(n298) );
  GTECH_XOR2 U281 ( .A(n312), .B(n275), .Z(n231) );
  GTECH_NOT U282 ( .A(n313), .Z(n275) );
  GTECH_OR_NOT U283 ( .A(n314), .B(I_b[7]), .Z(n313) );
  GTECH_OR_NOT U284 ( .A(n276), .B(I_b[6]), .Z(n312) );
  GTECH_NOT U285 ( .A(n270), .Z(n232) );
  GTECH_XOR3 U286 ( .A(n280), .B(n282), .C(n281), .Z(n270) );
  GTECH_OAI21 U287 ( .A(n315), .B(n316), .C(n317), .Z(n281) );
  GTECH_NOT U288 ( .A(n318), .Z(n282) );
  GTECH_OR_NOT U289 ( .A(n238), .B(I_b[5]), .Z(n318) );
  GTECH_NOT U290 ( .A(n278), .Z(n280) );
  GTECH_OR_NOT U291 ( .A(n200), .B(I_b[4]), .Z(n278) );
  GTECH_NOT U292 ( .A(n319), .Z(n272) );
  GTECH_NAND3 U293 ( .A(I_a[0]), .B(n320), .C(I_b[6]), .Z(n319) );
  GTECH_NOT U294 ( .A(n321), .Z(n320) );
  GTECH_XOR3 U295 ( .A(n265), .B(n266), .C(n294), .Z(n301) );
  GTECH_OAI21 U296 ( .A(n322), .B(n323), .C(n324), .Z(n294) );
  GTECH_OAI21 U297 ( .A(n325), .B(n326), .C(n327), .Z(n324) );
  GTECH_NOT U298 ( .A(n328), .Z(n266) );
  GTECH_OR_NOT U299 ( .A(n329), .B(I_a[6]), .Z(n328) );
  GTECH_NOT U300 ( .A(n292), .Z(n265) );
  GTECH_OR_NOT U301 ( .A(n330), .B(I_a[7]), .Z(n292) );
  GTECH_ADD_ABC U302 ( .A(n306), .B(n331), .C(n308), .COUT(n262) );
  GTECH_NOT U303 ( .A(n332), .Z(n308) );
  GTECH_XOR3 U304 ( .A(n325), .B(n327), .C(n322), .Z(n331) );
  GTECH_NOT U305 ( .A(n326), .Z(n322) );
  GTECH_XOR3 U306 ( .A(n287), .B(n289), .C(n288), .Z(n300) );
  GTECH_OAI21 U307 ( .A(n333), .B(n334), .C(n335), .Z(n288) );
  GTECH_OAI21 U308 ( .A(n336), .B(n337), .C(n338), .Z(n335) );
  GTECH_NOT U309 ( .A(n337), .Z(n333) );
  GTECH_NOT U310 ( .A(n339), .Z(n289) );
  GTECH_OR_NOT U311 ( .A(n176), .B(I_b[3]), .Z(n339) );
  GTECH_NOT U312 ( .A(n285), .Z(n287) );
  GTECH_OR_NOT U313 ( .A(n250), .B(I_a[5]), .Z(n285) );
  GTECH_NOT U314 ( .A(I_b[2]), .Z(n250) );
  GTECH_XOR2 U315 ( .A(n340), .B(n341), .Z(N146) );
  GTECH_XOR4 U316 ( .A(n307), .B(n332), .C(n305), .D(n306), .Z(n341) );
  GTECH_ADD_ABC U317 ( .A(n342), .B(n343), .C(n344), .COUT(n306) );
  GTECH_NOT U318 ( .A(n345), .Z(n344) );
  GTECH_XOR3 U319 ( .A(n346), .B(n347), .C(n348), .Z(n343) );
  GTECH_XOR2 U320 ( .A(n321), .B(n349), .Z(n305) );
  GTECH_AND2 U321 ( .A(I_b[6]), .B(I_a[0]), .Z(n349) );
  GTECH_XOR3 U322 ( .A(n350), .B(n351), .C(n317), .Z(n321) );
  GTECH_NAND3 U323 ( .A(I_b[4]), .B(I_a[1]), .C(n352), .Z(n317) );
  GTECH_NOT U324 ( .A(n316), .Z(n351) );
  GTECH_OR_NOT U325 ( .A(n276), .B(I_b[5]), .Z(n316) );
  GTECH_NOT U326 ( .A(n315), .Z(n350) );
  GTECH_OR_NOT U327 ( .A(n238), .B(I_b[4]), .Z(n315) );
  GTECH_XOR3 U328 ( .A(n336), .B(n338), .C(n337), .Z(n332) );
  GTECH_OAI21 U329 ( .A(n353), .B(n354), .C(n355), .Z(n337) );
  GTECH_OAI21 U330 ( .A(n356), .B(n357), .C(n358), .Z(n355) );
  GTECH_NOT U331 ( .A(n357), .Z(n353) );
  GTECH_NOT U332 ( .A(n359), .Z(n338) );
  GTECH_OR_NOT U333 ( .A(n200), .B(I_b[3]), .Z(n359) );
  GTECH_NOT U334 ( .A(n334), .Z(n336) );
  GTECH_OR_NOT U335 ( .A(n176), .B(I_b[2]), .Z(n334) );
  GTECH_NOT U336 ( .A(I_a[4]), .Z(n176) );
  GTECH_NOT U337 ( .A(n360), .Z(n307) );
  GTECH_XOR3 U338 ( .A(n325), .B(n327), .C(n326), .Z(n360) );
  GTECH_OAI21 U339 ( .A(n348), .B(n361), .C(n362), .Z(n326) );
  GTECH_OAI21 U340 ( .A(n346), .B(n363), .C(n347), .Z(n362) );
  GTECH_NOT U341 ( .A(n361), .Z(n346) );
  GTECH_NOT U342 ( .A(n363), .Z(n348) );
  GTECH_NOT U343 ( .A(n364), .Z(n327) );
  GTECH_OR_NOT U344 ( .A(n329), .B(I_a[5]), .Z(n364) );
  GTECH_NOT U345 ( .A(n323), .Z(n325) );
  GTECH_OR_NOT U346 ( .A(n330), .B(I_a[6]), .Z(n323) );
  GTECH_OA21 U347 ( .A(n309), .B(n310), .C(n311), .Z(n340) );
  GTECH_OAI21 U348 ( .A(n365), .B(n366), .C(n367), .Z(n311) );
  GTECH_NOT U349 ( .A(n309), .Z(n366) );
  GTECH_XOR3 U350 ( .A(n367), .B(n310), .C(n309), .Z(N145) );
  GTECH_XOR2 U351 ( .A(n368), .B(n352), .Z(n309) );
  GTECH_NOT U352 ( .A(n369), .Z(n352) );
  GTECH_OR_NOT U353 ( .A(n314), .B(I_b[5]), .Z(n369) );
  GTECH_OR_NOT U354 ( .A(n276), .B(I_b[4]), .Z(n368) );
  GTECH_NOT U355 ( .A(n365), .Z(n310) );
  GTECH_XOR2 U356 ( .A(n370), .B(n342), .Z(n365) );
  GTECH_ADD_ABC U357 ( .A(n371), .B(n372), .C(n373), .COUT(n342) );
  GTECH_XOR3 U358 ( .A(n374), .B(n375), .C(n376), .Z(n372) );
  GTECH_OA21 U359 ( .A(n377), .B(n378), .C(n379), .Z(n371) );
  GTECH_XOR4 U360 ( .A(n347), .B(n363), .C(n361), .D(n345), .Z(n370) );
  GTECH_XOR3 U361 ( .A(n356), .B(n358), .C(n357), .Z(n345) );
  GTECH_OAI21 U362 ( .A(n380), .B(n381), .C(n382), .Z(n357) );
  GTECH_NOT U363 ( .A(n383), .Z(n358) );
  GTECH_OR_NOT U364 ( .A(n238), .B(I_b[3]), .Z(n383) );
  GTECH_NOT U365 ( .A(n354), .Z(n356) );
  GTECH_OR_NOT U366 ( .A(n200), .B(I_b[2]), .Z(n354) );
  GTECH_OR_NOT U367 ( .A(n330), .B(I_a[5]), .Z(n361) );
  GTECH_OAI21 U368 ( .A(n376), .B(n384), .C(n385), .Z(n363) );
  GTECH_OAI21 U369 ( .A(n374), .B(n386), .C(n375), .Z(n385) );
  GTECH_NOT U370 ( .A(n386), .Z(n376) );
  GTECH_NOT U371 ( .A(n387), .Z(n347) );
  GTECH_OR_NOT U372 ( .A(n329), .B(I_a[4]), .Z(n387) );
  GTECH_NOT U373 ( .A(n388), .Z(n367) );
  GTECH_NAND3 U374 ( .A(I_a[0]), .B(n389), .C(I_b[4]), .Z(n388) );
  GTECH_XOR2 U375 ( .A(n390), .B(n389), .Z(N144) );
  GTECH_XOR2 U376 ( .A(n391), .B(n392), .Z(n389) );
  GTECH_XOR4 U377 ( .A(n375), .B(n386), .C(n373), .D(n374), .Z(n392) );
  GTECH_NOT U378 ( .A(n384), .Z(n374) );
  GTECH_OR_NOT U379 ( .A(n330), .B(I_a[4]), .Z(n384) );
  GTECH_NOT U380 ( .A(I_b[0]), .Z(n330) );
  GTECH_XOR3 U381 ( .A(n393), .B(n394), .C(n382), .Z(n373) );
  GTECH_NAND3 U382 ( .A(I_b[2]), .B(I_a[1]), .C(n395), .Z(n382) );
  GTECH_NOT U383 ( .A(n381), .Z(n394) );
  GTECH_OR_NOT U384 ( .A(n276), .B(I_b[3]), .Z(n381) );
  GTECH_NOT U385 ( .A(n380), .Z(n393) );
  GTECH_OR_NOT U386 ( .A(n238), .B(I_b[2]), .Z(n380) );
  GTECH_OAI21 U387 ( .A(n396), .B(n397), .C(n398), .Z(n386) );
  GTECH_OAI21 U388 ( .A(n399), .B(n400), .C(n401), .Z(n398) );
  GTECH_NOT U389 ( .A(n400), .Z(n396) );
  GTECH_NOT U390 ( .A(n402), .Z(n375) );
  GTECH_OR_NOT U391 ( .A(n329), .B(I_a[3]), .Z(n402) );
  GTECH_OA21 U392 ( .A(n377), .B(n378), .C(n379), .Z(n391) );
  GTECH_OAI21 U393 ( .A(n403), .B(n404), .C(n405), .Z(n379) );
  GTECH_NOT U394 ( .A(n377), .Z(n404) );
  GTECH_AND2 U395 ( .A(I_b[4]), .B(I_a[0]), .Z(n390) );
  GTECH_XOR3 U396 ( .A(n405), .B(n378), .C(n377), .Z(N143) );
  GTECH_XOR2 U397 ( .A(n406), .B(n395), .Z(n377) );
  GTECH_NOT U398 ( .A(n407), .Z(n395) );
  GTECH_OR_NOT U399 ( .A(n314), .B(I_b[3]), .Z(n407) );
  GTECH_NOT U400 ( .A(I_a[0]), .Z(n314) );
  GTECH_OR_NOT U401 ( .A(n276), .B(I_b[2]), .Z(n406) );
  GTECH_NOT U402 ( .A(I_a[1]), .Z(n276) );
  GTECH_NOT U403 ( .A(n403), .Z(n378) );
  GTECH_XOR3 U404 ( .A(n399), .B(n401), .C(n400), .Z(n403) );
  GTECH_OAI21 U405 ( .A(n408), .B(n409), .C(n410), .Z(n400) );
  GTECH_NOT U406 ( .A(n411), .Z(n401) );
  GTECH_OR_NOT U407 ( .A(n238), .B(I_b[1]), .Z(n411) );
  GTECH_NOT U408 ( .A(n397), .Z(n399) );
  GTECH_OR_NOT U409 ( .A(n200), .B(I_b[0]), .Z(n397) );
  GTECH_NOT U410 ( .A(I_a[3]), .Z(n200) );
  GTECH_NOT U411 ( .A(n412), .Z(n405) );
  GTECH_NAND3 U412 ( .A(I_a[0]), .B(n413), .C(I_b[2]), .Z(n412) );
  GTECH_XOR2 U413 ( .A(n414), .B(n413), .Z(N142) );
  GTECH_NOT U414 ( .A(n415), .Z(n413) );
  GTECH_XOR3 U415 ( .A(n416), .B(n417), .C(n410), .Z(n415) );
  GTECH_NAND3 U416 ( .A(n418), .B(I_b[0]), .C(I_a[1]), .Z(n410) );
  GTECH_NOT U417 ( .A(n408), .Z(n417) );
  GTECH_OR_NOT U418 ( .A(n329), .B(I_a[1]), .Z(n408) );
  GTECH_NOT U419 ( .A(n409), .Z(n416) );
  GTECH_OR_NOT U420 ( .A(n238), .B(I_b[0]), .Z(n409) );
  GTECH_NOT U421 ( .A(I_a[2]), .Z(n238) );
  GTECH_AND2 U422 ( .A(I_b[2]), .B(I_a[0]), .Z(n414) );
  GTECH_XOR2 U423 ( .A(n418), .B(n419), .Z(N141) );
  GTECH_AND2 U424 ( .A(I_a[1]), .B(I_b[0]), .Z(n419) );
  GTECH_NOT U425 ( .A(n420), .Z(n418) );
  GTECH_OR_NOT U426 ( .A(n329), .B(I_a[0]), .Z(n420) );
  GTECH_NOT U427 ( .A(I_b[1]), .Z(n329) );
  GTECH_AND2 U428 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

