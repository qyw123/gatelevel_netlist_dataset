
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n85) );
  GTECH_XNOR2 U78 ( .A(n84), .B(n90), .Z(N154) );
  GTECH_XNOR2 U79 ( .A(n91), .B(n92), .Z(n90) );
  GTECH_NOT U80 ( .A(n86), .Z(n92) );
  GTECH_XNOR2 U81 ( .A(n93), .B(n88), .Z(n86) );
  GTECH_NOT U82 ( .A(n94), .Z(n88) );
  GTECH_OR_NOT U83 ( .A(n95), .B(I_b[7]), .Z(n94) );
  GTECH_NOT U84 ( .A(n89), .Z(n93) );
  GTECH_OAI21 U85 ( .A(n96), .B(n97), .C(n98), .Z(n89) );
  GTECH_OAI21 U86 ( .A(n99), .B(n100), .C(n101), .Z(n98) );
  GTECH_NOT U87 ( .A(n100), .Z(n96) );
  GTECH_NOT U88 ( .A(n87), .Z(n91) );
  GTECH_OAI2N2 U89 ( .A(n102), .B(n103), .C(n104), .D(n105), .Z(n87) );
  GTECH_OR_NOT U90 ( .A(n106), .B(n102), .Z(n105) );
  GTECH_NOT U91 ( .A(n107), .Z(n84) );
  GTECH_OR_NOT U92 ( .A(n108), .B(n109), .Z(n107) );
  GTECH_NOT U93 ( .A(n110), .Z(n109) );
  GTECH_XNOR2 U94 ( .A(n111), .B(n110), .Z(N153) );
  GTECH_XOR3 U95 ( .A(n106), .B(n102), .C(n104), .Z(n110) );
  GTECH_XOR3 U96 ( .A(n99), .B(n101), .C(n100), .Z(n104) );
  GTECH_OAI21 U97 ( .A(n112), .B(n113), .C(n114), .Z(n100) );
  GTECH_OAI21 U98 ( .A(n115), .B(n116), .C(n117), .Z(n114) );
  GTECH_NOT U99 ( .A(n116), .Z(n112) );
  GTECH_NOT U100 ( .A(n118), .Z(n101) );
  GTECH_OR_NOT U101 ( .A(n119), .B(I_b[7]), .Z(n118) );
  GTECH_NOT U102 ( .A(n97), .Z(n99) );
  GTECH_OR_NOT U103 ( .A(n120), .B(I_a[7]), .Z(n97) );
  GTECH_NOT U104 ( .A(I_b[6]), .Z(n120) );
  GTECH_ADD_ABC U105 ( .A(n121), .B(n122), .C(n123), .COUT(n102) );
  GTECH_NOT U106 ( .A(n124), .Z(n123) );
  GTECH_XNOR2 U107 ( .A(n125), .B(n126), .Z(n122) );
  GTECH_OR_NOT U108 ( .A(n127), .B(I_a[7]), .Z(n126) );
  GTECH_NOT U109 ( .A(n103), .Z(n106) );
  GTECH_OR_NOT U110 ( .A(n125), .B(I_a[7]), .Z(n103) );
  GTECH_NOT U111 ( .A(n108), .Z(n111) );
  GTECH_OR_NOT U112 ( .A(n128), .B(n129), .Z(n108) );
  GTECH_XNOR2 U113 ( .A(n128), .B(n129), .Z(N152) );
  GTECH_XOR4 U114 ( .A(n125), .B(n130), .C(n121), .D(n124), .Z(n129) );
  GTECH_XOR3 U115 ( .A(n115), .B(n117), .C(n116), .Z(n124) );
  GTECH_OAI21 U116 ( .A(n131), .B(n132), .C(n133), .Z(n116) );
  GTECH_OAI21 U117 ( .A(n134), .B(n135), .C(n136), .Z(n133) );
  GTECH_NOT U118 ( .A(n135), .Z(n131) );
  GTECH_NOT U119 ( .A(n137), .Z(n117) );
  GTECH_OR_NOT U120 ( .A(n138), .B(I_b[7]), .Z(n137) );
  GTECH_NOT U121 ( .A(n113), .Z(n115) );
  GTECH_OR_NOT U122 ( .A(n119), .B(I_b[6]), .Z(n113) );
  GTECH_NOT U123 ( .A(I_a[6]), .Z(n119) );
  GTECH_ADD_ABC U124 ( .A(n139), .B(n140), .C(n141), .COUT(n121) );
  GTECH_NOT U125 ( .A(n142), .Z(n141) );
  GTECH_XOR3 U126 ( .A(n143), .B(n144), .C(n145), .Z(n140) );
  GTECH_AND2 U127 ( .A(I_a[7]), .B(I_b[5]), .Z(n130) );
  GTECH_OA21 U128 ( .A(n145), .B(n146), .C(n147), .Z(n125) );
  GTECH_OAI21 U129 ( .A(n143), .B(n148), .C(n144), .Z(n147) );
  GTECH_NOT U130 ( .A(n146), .Z(n143) );
  GTECH_NOT U131 ( .A(n148), .Z(n145) );
  GTECH_ADD_ABC U132 ( .A(n149), .B(n150), .C(n151), .COUT(n128) );
  GTECH_NOT U133 ( .A(n152), .Z(n151) );
  GTECH_OA22 U134 ( .A(n153), .B(n95), .C(n154), .D(n155), .Z(n150) );
  GTECH_OA21 U135 ( .A(n156), .B(n157), .C(n158), .Z(n149) );
  GTECH_XOR3 U136 ( .A(n159), .B(n152), .C(n160), .Z(N151) );
  GTECH_OA21 U137 ( .A(n156), .B(n157), .C(n158), .Z(n160) );
  GTECH_OAI21 U138 ( .A(n161), .B(n162), .C(n163), .Z(n158) );
  GTECH_XOR3 U139 ( .A(n142), .B(n139), .C(n164), .Z(n152) );
  GTECH_XOR3 U140 ( .A(n144), .B(n148), .C(n146), .Z(n164) );
  GTECH_OR_NOT U141 ( .A(n165), .B(I_a[7]), .Z(n146) );
  GTECH_OAI21 U142 ( .A(n166), .B(n167), .C(n168), .Z(n148) );
  GTECH_OAI21 U143 ( .A(n169), .B(n170), .C(n171), .Z(n168) );
  GTECH_NOT U144 ( .A(n172), .Z(n144) );
  GTECH_OR_NOT U145 ( .A(n127), .B(I_a[6]), .Z(n172) );
  GTECH_ADD_ABC U146 ( .A(n173), .B(n174), .C(n175), .COUT(n139) );
  GTECH_NOT U147 ( .A(n176), .Z(n175) );
  GTECH_XOR3 U148 ( .A(n169), .B(n171), .C(n166), .Z(n174) );
  GTECH_NOT U149 ( .A(n170), .Z(n166) );
  GTECH_NOT U150 ( .A(n167), .Z(n169) );
  GTECH_XOR3 U151 ( .A(n134), .B(n136), .C(n135), .Z(n142) );
  GTECH_OAI21 U152 ( .A(n177), .B(n178), .C(n179), .Z(n135) );
  GTECH_OAI21 U153 ( .A(n180), .B(n181), .C(n182), .Z(n179) );
  GTECH_NOT U154 ( .A(n181), .Z(n177) );
  GTECH_NOT U155 ( .A(n183), .Z(n136) );
  GTECH_OR_NOT U156 ( .A(n184), .B(I_b[7]), .Z(n183) );
  GTECH_NOT U157 ( .A(n132), .Z(n134) );
  GTECH_OR_NOT U158 ( .A(n138), .B(I_b[6]), .Z(n132) );
  GTECH_NOT U159 ( .A(I_a[5]), .Z(n138) );
  GTECH_OA22 U160 ( .A(n153), .B(n95), .C(n154), .D(n155), .Z(n159) );
  GTECH_NOT U161 ( .A(I_a[7]), .Z(n95) );
  GTECH_XOR3 U162 ( .A(n156), .B(n161), .C(n185), .Z(N150) );
  GTECH_NOT U163 ( .A(n163), .Z(n185) );
  GTECH_XOR3 U164 ( .A(n176), .B(n173), .C(n186), .Z(n163) );
  GTECH_XOR3 U165 ( .A(n171), .B(n170), .C(n167), .Z(n186) );
  GTECH_OR_NOT U166 ( .A(n165), .B(I_a[6]), .Z(n167) );
  GTECH_OAI21 U167 ( .A(n187), .B(n188), .C(n189), .Z(n170) );
  GTECH_OAI21 U168 ( .A(n190), .B(n191), .C(n192), .Z(n189) );
  GTECH_NOT U169 ( .A(n193), .Z(n171) );
  GTECH_OR_NOT U170 ( .A(n127), .B(I_a[5]), .Z(n193) );
  GTECH_NOT U171 ( .A(I_b[5]), .Z(n127) );
  GTECH_ADD_ABC U172 ( .A(n194), .B(n195), .C(n196), .COUT(n173) );
  GTECH_NOT U173 ( .A(n197), .Z(n196) );
  GTECH_XOR3 U174 ( .A(n190), .B(n192), .C(n187), .Z(n195) );
  GTECH_NOT U175 ( .A(n191), .Z(n187) );
  GTECH_NOT U176 ( .A(n188), .Z(n190) );
  GTECH_XOR3 U177 ( .A(n180), .B(n182), .C(n181), .Z(n176) );
  GTECH_OAI21 U178 ( .A(n198), .B(n199), .C(n200), .Z(n181) );
  GTECH_OAI21 U179 ( .A(n201), .B(n202), .C(n203), .Z(n200) );
  GTECH_NOT U180 ( .A(n202), .Z(n198) );
  GTECH_NOT U181 ( .A(n204), .Z(n182) );
  GTECH_OR_NOT U182 ( .A(n205), .B(I_b[7]), .Z(n204) );
  GTECH_NOT U183 ( .A(n178), .Z(n180) );
  GTECH_OR_NOT U184 ( .A(n184), .B(I_b[6]), .Z(n178) );
  GTECH_NOT U185 ( .A(n157), .Z(n161) );
  GTECH_XNOR2 U186 ( .A(n154), .B(n155), .Z(n157) );
  GTECH_ADD_AB U187 ( .A(n153), .B(n206), .S(n155) );
  GTECH_AND2 U188 ( .A(I_a[7]), .B(I_b[3]), .Z(n206) );
  GTECH_AND2 U189 ( .A(n207), .B(n208), .Z(n153) );
  GTECH_OR_NOT U190 ( .A(n209), .B(n210), .Z(n208) );
  GTECH_OAI21 U191 ( .A(n211), .B(n210), .C(n212), .Z(n207) );
  GTECH_AOI2N2 U192 ( .A(n213), .B(n214), .C(n215), .D(n216), .Z(n154) );
  GTECH_OR_NOT U193 ( .A(n217), .B(n215), .Z(n214) );
  GTECH_NOT U194 ( .A(n162), .Z(n156) );
  GTECH_OAI2N2 U195 ( .A(n218), .B(n219), .C(n220), .D(n221), .Z(n162) );
  GTECH_OR_NOT U196 ( .A(n222), .B(n218), .Z(n221) );
  GTECH_XOR3 U197 ( .A(n218), .B(n222), .C(n223), .Z(N149) );
  GTECH_NOT U198 ( .A(n220), .Z(n223) );
  GTECH_XOR3 U199 ( .A(n197), .B(n194), .C(n224), .Z(n220) );
  GTECH_XOR3 U200 ( .A(n192), .B(n191), .C(n188), .Z(n224) );
  GTECH_OR_NOT U201 ( .A(n165), .B(I_a[5]), .Z(n188) );
  GTECH_NOT U202 ( .A(I_b[4]), .Z(n165) );
  GTECH_OAI21 U203 ( .A(n225), .B(n226), .C(n227), .Z(n191) );
  GTECH_OAI21 U204 ( .A(n228), .B(n229), .C(n230), .Z(n227) );
  GTECH_NOT U205 ( .A(n231), .Z(n192) );
  GTECH_OR_NOT U206 ( .A(n184), .B(I_b[5]), .Z(n231) );
  GTECH_ADD_ABC U207 ( .A(n232), .B(n233), .C(n234), .COUT(n194) );
  GTECH_XOR3 U208 ( .A(n228), .B(n230), .C(n225), .Z(n233) );
  GTECH_NOT U209 ( .A(n229), .Z(n225) );
  GTECH_OA21 U210 ( .A(n235), .B(n236), .C(n237), .Z(n232) );
  GTECH_XOR3 U211 ( .A(n201), .B(n203), .C(n202), .Z(n197) );
  GTECH_OAI21 U212 ( .A(n238), .B(n239), .C(n240), .Z(n202) );
  GTECH_NOT U213 ( .A(n241), .Z(n203) );
  GTECH_OR_NOT U214 ( .A(n242), .B(I_b[7]), .Z(n241) );
  GTECH_NOT U215 ( .A(n199), .Z(n201) );
  GTECH_OR_NOT U216 ( .A(n205), .B(I_b[6]), .Z(n199) );
  GTECH_NOT U217 ( .A(n219), .Z(n222) );
  GTECH_XOR3 U218 ( .A(n217), .B(n215), .C(n213), .Z(n219) );
  GTECH_XOR3 U219 ( .A(n211), .B(n212), .C(n210), .Z(n213) );
  GTECH_OAI21 U220 ( .A(n243), .B(n244), .C(n245), .Z(n210) );
  GTECH_OAI21 U221 ( .A(n246), .B(n247), .C(n248), .Z(n245) );
  GTECH_NOT U222 ( .A(n247), .Z(n243) );
  GTECH_NOT U223 ( .A(n249), .Z(n212) );
  GTECH_OR_NOT U224 ( .A(n250), .B(I_a[6]), .Z(n249) );
  GTECH_NOT U225 ( .A(n209), .Z(n211) );
  GTECH_OR_NOT U226 ( .A(n251), .B(I_a[7]), .Z(n209) );
  GTECH_ADD_ABC U227 ( .A(n252), .B(n253), .C(n254), .COUT(n215) );
  GTECH_XNOR2 U228 ( .A(n255), .B(n256), .Z(n253) );
  GTECH_OR_NOT U229 ( .A(n257), .B(I_a[7]), .Z(n256) );
  GTECH_NOT U230 ( .A(n216), .Z(n217) );
  GTECH_OR_NOT U231 ( .A(n255), .B(I_a[7]), .Z(n216) );
  GTECH_ADD_ABC U232 ( .A(n258), .B(n259), .C(n260), .COUT(n218) );
  GTECH_XOR3 U233 ( .A(n252), .B(n261), .C(n254), .Z(n259) );
  GTECH_NOT U234 ( .A(n262), .Z(n254) );
  GTECH_XOR3 U235 ( .A(n263), .B(n260), .C(n258), .Z(N148) );
  GTECH_ADD_ABC U236 ( .A(n264), .B(n265), .C(n266), .COUT(n258) );
  GTECH_NOT U237 ( .A(n267), .Z(n266) );
  GTECH_XOR3 U238 ( .A(n268), .B(n269), .C(n270), .Z(n265) );
  GTECH_NOT U239 ( .A(n271), .Z(n269) );
  GTECH_XOR3 U240 ( .A(n272), .B(n234), .C(n273), .Z(n260) );
  GTECH_OAI21 U241 ( .A(n235), .B(n236), .C(n237), .Z(n273) );
  GTECH_OAI21 U242 ( .A(n274), .B(n275), .C(n276), .Z(n237) );
  GTECH_NOT U243 ( .A(n235), .Z(n275) );
  GTECH_XOR3 U244 ( .A(n277), .B(n278), .C(n240), .Z(n234) );
  GTECH_NAND3 U245 ( .A(I_b[6]), .B(I_a[1]), .C(n279), .Z(n240) );
  GTECH_NOT U246 ( .A(n239), .Z(n278) );
  GTECH_OR_NOT U247 ( .A(n280), .B(I_b[7]), .Z(n239) );
  GTECH_NOT U248 ( .A(n238), .Z(n277) );
  GTECH_OR_NOT U249 ( .A(n242), .B(I_b[6]), .Z(n238) );
  GTECH_XOR3 U250 ( .A(n230), .B(n229), .C(n228), .Z(n272) );
  GTECH_NOT U251 ( .A(n226), .Z(n228) );
  GTECH_OR_NOT U252 ( .A(n184), .B(I_b[4]), .Z(n226) );
  GTECH_OAI21 U253 ( .A(n281), .B(n282), .C(n283), .Z(n229) );
  GTECH_OAI21 U254 ( .A(n284), .B(n285), .C(n286), .Z(n283) );
  GTECH_NOT U255 ( .A(n285), .Z(n281) );
  GTECH_NOT U256 ( .A(n287), .Z(n230) );
  GTECH_OR_NOT U257 ( .A(n205), .B(I_b[5]), .Z(n287) );
  GTECH_XOR3 U258 ( .A(n261), .B(n262), .C(n252), .Z(n263) );
  GTECH_ADD_ABC U259 ( .A(n268), .B(n288), .C(n270), .COUT(n252) );
  GTECH_NOT U260 ( .A(n289), .Z(n270) );
  GTECH_XOR3 U261 ( .A(n290), .B(n291), .C(n292), .Z(n288) );
  GTECH_XOR3 U262 ( .A(n246), .B(n248), .C(n247), .Z(n262) );
  GTECH_OAI21 U263 ( .A(n293), .B(n294), .C(n295), .Z(n247) );
  GTECH_OAI21 U264 ( .A(n296), .B(n297), .C(n298), .Z(n295) );
  GTECH_NOT U265 ( .A(n297), .Z(n293) );
  GTECH_NOT U266 ( .A(n299), .Z(n248) );
  GTECH_OR_NOT U267 ( .A(n250), .B(I_a[5]), .Z(n299) );
  GTECH_NOT U268 ( .A(I_b[3]), .Z(n250) );
  GTECH_NOT U269 ( .A(n244), .Z(n246) );
  GTECH_OR_NOT U270 ( .A(n251), .B(I_a[6]), .Z(n244) );
  GTECH_ADD_AB U271 ( .A(n255), .B(n300), .S(n261) );
  GTECH_AND2 U272 ( .A(I_a[7]), .B(I_b[1]), .Z(n300) );
  GTECH_OA21 U273 ( .A(n292), .B(n301), .C(n302), .Z(n255) );
  GTECH_OAI21 U274 ( .A(n290), .B(n303), .C(n291), .Z(n302) );
  GTECH_NOT U275 ( .A(n303), .Z(n292) );
  GTECH_XOR3 U276 ( .A(n267), .B(n264), .C(n304), .Z(N147) );
  GTECH_XOR3 U277 ( .A(n289), .B(n268), .C(n271), .Z(n304) );
  GTECH_XOR3 U278 ( .A(n290), .B(n291), .C(n303), .Z(n271) );
  GTECH_OAI21 U279 ( .A(n305), .B(n306), .C(n307), .Z(n303) );
  GTECH_OAI21 U280 ( .A(n308), .B(n309), .C(n310), .Z(n307) );
  GTECH_NOT U281 ( .A(n311), .Z(n291) );
  GTECH_OR_NOT U282 ( .A(n257), .B(I_a[6]), .Z(n311) );
  GTECH_NOT U283 ( .A(n301), .Z(n290) );
  GTECH_OR_NOT U284 ( .A(n312), .B(I_a[7]), .Z(n301) );
  GTECH_ADD_ABC U285 ( .A(n313), .B(n314), .C(n315), .COUT(n268) );
  GTECH_XOR3 U286 ( .A(n308), .B(n310), .C(n305), .Z(n314) );
  GTECH_NOT U287 ( .A(n309), .Z(n305) );
  GTECH_XOR3 U288 ( .A(n296), .B(n298), .C(n297), .Z(n289) );
  GTECH_OAI21 U289 ( .A(n316), .B(n317), .C(n318), .Z(n297) );
  GTECH_OAI21 U290 ( .A(n319), .B(n320), .C(n321), .Z(n318) );
  GTECH_NOT U291 ( .A(n320), .Z(n316) );
  GTECH_NOT U292 ( .A(n322), .Z(n298) );
  GTECH_OR_NOT U293 ( .A(n184), .B(I_b[3]), .Z(n322) );
  GTECH_NOT U294 ( .A(n294), .Z(n296) );
  GTECH_OR_NOT U295 ( .A(n251), .B(I_a[5]), .Z(n294) );
  GTECH_NOT U296 ( .A(I_b[2]), .Z(n251) );
  GTECH_ADD_ABC U297 ( .A(n323), .B(n324), .C(n325), .COUT(n264) );
  GTECH_XOR3 U298 ( .A(n313), .B(n326), .C(n315), .Z(n324) );
  GTECH_NOT U299 ( .A(n327), .Z(n315) );
  GTECH_OA21 U300 ( .A(n328), .B(n329), .C(n330), .Z(n323) );
  GTECH_XOR3 U301 ( .A(n276), .B(n236), .C(n235), .Z(n267) );
  GTECH_XNOR2 U302 ( .A(n279), .B(n331), .Z(n235) );
  GTECH_AND2 U303 ( .A(I_b[6]), .B(I_a[1]), .Z(n331) );
  GTECH_NOT U304 ( .A(n332), .Z(n279) );
  GTECH_OR_NOT U305 ( .A(n333), .B(I_b[7]), .Z(n332) );
  GTECH_NOT U306 ( .A(n274), .Z(n236) );
  GTECH_XOR3 U307 ( .A(n284), .B(n286), .C(n285), .Z(n274) );
  GTECH_OAI21 U308 ( .A(n334), .B(n335), .C(n336), .Z(n285) );
  GTECH_NOT U309 ( .A(n337), .Z(n286) );
  GTECH_OR_NOT U310 ( .A(n242), .B(I_b[5]), .Z(n337) );
  GTECH_NOT U311 ( .A(n282), .Z(n284) );
  GTECH_OR_NOT U312 ( .A(n205), .B(I_b[4]), .Z(n282) );
  GTECH_NOT U313 ( .A(n338), .Z(n276) );
  GTECH_NAND3 U314 ( .A(I_a[0]), .B(n339), .C(I_b[6]), .Z(n338) );
  GTECH_XOR3 U315 ( .A(n340), .B(n325), .C(n341), .Z(N146) );
  GTECH_OA21 U316 ( .A(n328), .B(n329), .C(n330), .Z(n341) );
  GTECH_OAI21 U317 ( .A(n342), .B(n343), .C(n344), .Z(n330) );
  GTECH_NOT U318 ( .A(n328), .Z(n343) );
  GTECH_XNOR2 U319 ( .A(n345), .B(n339), .Z(n325) );
  GTECH_NOT U320 ( .A(n346), .Z(n339) );
  GTECH_XOR3 U321 ( .A(n347), .B(n348), .C(n336), .Z(n346) );
  GTECH_NAND3 U322 ( .A(I_b[4]), .B(I_a[1]), .C(n349), .Z(n336) );
  GTECH_NOT U323 ( .A(n335), .Z(n348) );
  GTECH_OR_NOT U324 ( .A(n280), .B(I_b[5]), .Z(n335) );
  GTECH_NOT U325 ( .A(n334), .Z(n347) );
  GTECH_OR_NOT U326 ( .A(n242), .B(I_b[4]), .Z(n334) );
  GTECH_AND2 U327 ( .A(I_b[6]), .B(I_a[0]), .Z(n345) );
  GTECH_XOR3 U328 ( .A(n326), .B(n327), .C(n313), .Z(n340) );
  GTECH_ADD_ABC U329 ( .A(n350), .B(n351), .C(n352), .COUT(n313) );
  GTECH_NOT U330 ( .A(n353), .Z(n352) );
  GTECH_XOR3 U331 ( .A(n354), .B(n355), .C(n356), .Z(n351) );
  GTECH_XOR3 U332 ( .A(n319), .B(n321), .C(n320), .Z(n327) );
  GTECH_OAI21 U333 ( .A(n357), .B(n358), .C(n359), .Z(n320) );
  GTECH_OAI21 U334 ( .A(n360), .B(n361), .C(n362), .Z(n359) );
  GTECH_NOT U335 ( .A(n361), .Z(n357) );
  GTECH_NOT U336 ( .A(n363), .Z(n321) );
  GTECH_OR_NOT U337 ( .A(n205), .B(I_b[3]), .Z(n363) );
  GTECH_NOT U338 ( .A(n317), .Z(n319) );
  GTECH_OR_NOT U339 ( .A(n184), .B(I_b[2]), .Z(n317) );
  GTECH_NOT U340 ( .A(I_a[4]), .Z(n184) );
  GTECH_NOT U341 ( .A(n364), .Z(n326) );
  GTECH_XOR3 U342 ( .A(n308), .B(n310), .C(n309), .Z(n364) );
  GTECH_OAI21 U343 ( .A(n356), .B(n365), .C(n366), .Z(n309) );
  GTECH_OAI21 U344 ( .A(n354), .B(n367), .C(n355), .Z(n366) );
  GTECH_NOT U345 ( .A(n365), .Z(n354) );
  GTECH_NOT U346 ( .A(n367), .Z(n356) );
  GTECH_NOT U347 ( .A(n368), .Z(n310) );
  GTECH_OR_NOT U348 ( .A(n257), .B(I_a[5]), .Z(n368) );
  GTECH_NOT U349 ( .A(n306), .Z(n308) );
  GTECH_OR_NOT U350 ( .A(n312), .B(I_a[6]), .Z(n306) );
  GTECH_XOR3 U351 ( .A(n344), .B(n329), .C(n328), .Z(N145) );
  GTECH_XNOR2 U352 ( .A(n349), .B(n369), .Z(n328) );
  GTECH_AND2 U353 ( .A(I_b[4]), .B(I_a[1]), .Z(n369) );
  GTECH_NOT U354 ( .A(n370), .Z(n349) );
  GTECH_OR_NOT U355 ( .A(n333), .B(I_b[5]), .Z(n370) );
  GTECH_NOT U356 ( .A(n342), .Z(n329) );
  GTECH_XOR3 U357 ( .A(n353), .B(n350), .C(n371), .Z(n342) );
  GTECH_XOR3 U358 ( .A(n355), .B(n367), .C(n365), .Z(n371) );
  GTECH_OR_NOT U359 ( .A(n312), .B(I_a[5]), .Z(n365) );
  GTECH_OAI21 U360 ( .A(n372), .B(n373), .C(n374), .Z(n367) );
  GTECH_OAI21 U361 ( .A(n375), .B(n376), .C(n377), .Z(n374) );
  GTECH_NOT U362 ( .A(n378), .Z(n355) );
  GTECH_OR_NOT U363 ( .A(n257), .B(I_a[4]), .Z(n378) );
  GTECH_ADD_ABC U364 ( .A(n379), .B(n380), .C(n381), .COUT(n350) );
  GTECH_XOR3 U365 ( .A(n375), .B(n377), .C(n372), .Z(n380) );
  GTECH_NOT U366 ( .A(n376), .Z(n372) );
  GTECH_OA21 U367 ( .A(n382), .B(n383), .C(n384), .Z(n379) );
  GTECH_XOR3 U368 ( .A(n360), .B(n362), .C(n361), .Z(n353) );
  GTECH_OAI21 U369 ( .A(n385), .B(n386), .C(n387), .Z(n361) );
  GTECH_NOT U370 ( .A(n388), .Z(n362) );
  GTECH_OR_NOT U371 ( .A(n242), .B(I_b[3]), .Z(n388) );
  GTECH_NOT U372 ( .A(n358), .Z(n360) );
  GTECH_OR_NOT U373 ( .A(n205), .B(I_b[2]), .Z(n358) );
  GTECH_NOT U374 ( .A(n389), .Z(n344) );
  GTECH_NAND3 U375 ( .A(I_a[0]), .B(n390), .C(I_b[4]), .Z(n389) );
  GTECH_NOT U376 ( .A(n391), .Z(n390) );
  GTECH_XNOR2 U377 ( .A(n392), .B(n391), .Z(N144) );
  GTECH_XOR3 U378 ( .A(n393), .B(n381), .C(n394), .Z(n391) );
  GTECH_OAI21 U379 ( .A(n382), .B(n383), .C(n384), .Z(n394) );
  GTECH_OAI21 U380 ( .A(n395), .B(n396), .C(n397), .Z(n384) );
  GTECH_NOT U381 ( .A(n382), .Z(n396) );
  GTECH_XOR3 U382 ( .A(n398), .B(n399), .C(n387), .Z(n381) );
  GTECH_NAND3 U383 ( .A(I_b[2]), .B(I_a[1]), .C(n400), .Z(n387) );
  GTECH_NOT U384 ( .A(n386), .Z(n399) );
  GTECH_OR_NOT U385 ( .A(n280), .B(I_b[3]), .Z(n386) );
  GTECH_NOT U386 ( .A(I_a[1]), .Z(n280) );
  GTECH_NOT U387 ( .A(n385), .Z(n398) );
  GTECH_OR_NOT U388 ( .A(n242), .B(I_b[2]), .Z(n385) );
  GTECH_XOR3 U389 ( .A(n377), .B(n376), .C(n375), .Z(n393) );
  GTECH_NOT U390 ( .A(n373), .Z(n375) );
  GTECH_OR_NOT U391 ( .A(n312), .B(I_a[4]), .Z(n373) );
  GTECH_OAI21 U392 ( .A(n401), .B(n402), .C(n403), .Z(n376) );
  GTECH_OAI21 U393 ( .A(n404), .B(n405), .C(n406), .Z(n403) );
  GTECH_NOT U394 ( .A(n405), .Z(n401) );
  GTECH_NOT U395 ( .A(n407), .Z(n377) );
  GTECH_OR_NOT U396 ( .A(n257), .B(I_a[3]), .Z(n407) );
  GTECH_AND2 U397 ( .A(I_b[4]), .B(I_a[0]), .Z(n392) );
  GTECH_XOR3 U398 ( .A(n397), .B(n383), .C(n382), .Z(N143) );
  GTECH_XNOR2 U399 ( .A(n400), .B(n408), .Z(n382) );
  GTECH_AND2 U400 ( .A(I_b[2]), .B(I_a[1]), .Z(n408) );
  GTECH_NOT U401 ( .A(n409), .Z(n400) );
  GTECH_OR_NOT U402 ( .A(n333), .B(I_b[3]), .Z(n409) );
  GTECH_NOT U403 ( .A(I_a[0]), .Z(n333) );
  GTECH_NOT U404 ( .A(n395), .Z(n383) );
  GTECH_XOR3 U405 ( .A(n404), .B(n406), .C(n405), .Z(n395) );
  GTECH_OAI21 U406 ( .A(n410), .B(n411), .C(n412), .Z(n405) );
  GTECH_NOT U407 ( .A(n413), .Z(n406) );
  GTECH_OR_NOT U408 ( .A(n242), .B(I_b[1]), .Z(n413) );
  GTECH_NOT U409 ( .A(n402), .Z(n404) );
  GTECH_OR_NOT U410 ( .A(n205), .B(I_b[0]), .Z(n402) );
  GTECH_NOT U411 ( .A(I_a[3]), .Z(n205) );
  GTECH_NOT U412 ( .A(n414), .Z(n397) );
  GTECH_NAND3 U413 ( .A(I_a[0]), .B(n415), .C(I_b[2]), .Z(n414) );
  GTECH_NOT U414 ( .A(n416), .Z(n415) );
  GTECH_XNOR2 U415 ( .A(n417), .B(n416), .Z(N142) );
  GTECH_XOR3 U416 ( .A(n418), .B(n419), .C(n412), .Z(n416) );
  GTECH_NAND3 U417 ( .A(n420), .B(I_b[0]), .C(I_a[1]), .Z(n412) );
  GTECH_NOT U418 ( .A(n410), .Z(n419) );
  GTECH_OR_NOT U419 ( .A(n257), .B(I_a[1]), .Z(n410) );
  GTECH_NOT U420 ( .A(n411), .Z(n418) );
  GTECH_OR_NOT U421 ( .A(n242), .B(I_b[0]), .Z(n411) );
  GTECH_NOT U422 ( .A(I_a[2]), .Z(n242) );
  GTECH_AND2 U423 ( .A(I_b[2]), .B(I_a[0]), .Z(n417) );
  GTECH_XNOR2 U424 ( .A(n420), .B(n421), .Z(N141) );
  GTECH_OR_NOT U425 ( .A(n312), .B(I_a[1]), .Z(n421) );
  GTECH_NOT U426 ( .A(I_b[0]), .Z(n312) );
  GTECH_NOT U427 ( .A(n422), .Z(n420) );
  GTECH_OR_NOT U428 ( .A(n257), .B(I_a[0]), .Z(n422) );
  GTECH_NOT U429 ( .A(I_b[1]), .Z(n257) );
  GTECH_AND2 U430 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

