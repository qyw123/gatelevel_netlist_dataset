
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383;

  GTECH_MUX2 U129 ( .A(n268), .B(n269), .S(n270), .Z(sum[9]) );
  GTECH_XOR2 U130 ( .A(n271), .B(n272), .Z(n269) );
  GTECH_XOR2 U131 ( .A(n273), .B(n271), .Z(n268) );
  GTECH_OR_NOT U132 ( .A(n274), .B(n275), .Z(n271) );
  GTECH_XNOR2 U133 ( .A(n270), .B(n276), .Z(sum[8]) );
  GTECH_MUX2 U134 ( .A(n277), .B(n278), .S(n279), .Z(sum[7]) );
  GTECH_XOR2 U135 ( .A(n280), .B(n281), .Z(n278) );
  GTECH_AOI21 U136 ( .A(n282), .B(n283), .C(n284), .Z(n280) );
  GTECH_OA21 U137 ( .A(n283), .B(n282), .C(n285), .Z(n284) );
  GTECH_XNOR2 U138 ( .A(n281), .B(n286), .Z(n277) );
  GTECH_XOR2 U139 ( .A(a[7]), .B(b[7]), .Z(n281) );
  GTECH_XNOR3 U140 ( .A(n285), .B(a[6]), .C(n287), .Z(sum[6]) );
  GTECH_OAI21 U141 ( .A(n279), .B(n288), .C(n283), .Z(n287) );
  GTECH_AOI21 U142 ( .A(n289), .B(n290), .C(n291), .Z(n283) );
  GTECH_NOT U143 ( .A(b[6]), .Z(n285) );
  GTECH_MUX2 U144 ( .A(n292), .B(n293), .S(n294), .Z(sum[5]) );
  GTECH_OR_NOT U145 ( .A(n291), .B(n289), .Z(n294) );
  GTECH_NOT U146 ( .A(n295), .Z(n293) );
  GTECH_AOI21 U147 ( .A(n296), .B(n297), .C(n290), .Z(n295) );
  GTECH_NOR2 U148 ( .A(n298), .B(n299), .Z(n290) );
  GTECH_OAI21 U149 ( .A(a[4]), .B(n296), .C(n300), .Z(n292) );
  GTECH_OAI21 U150 ( .A(n279), .B(n298), .C(n299), .Z(n300) );
  GTECH_XOR2 U151 ( .A(n301), .B(n296), .Z(sum[4]) );
  GTECH_MUX2 U152 ( .A(n302), .B(n303), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U153 ( .A(n304), .B(n305), .Z(n303) );
  GTECH_XNOR2 U154 ( .A(n306), .B(n304), .Z(n302) );
  GTECH_XNOR2 U155 ( .A(a[3]), .B(b[3]), .Z(n304) );
  GTECH_AOI21 U156 ( .A(n307), .B(n308), .C(n309), .Z(n306) );
  GTECH_OA21 U157 ( .A(n308), .B(n307), .C(n310), .Z(n309) );
  GTECH_MUX2 U158 ( .A(n311), .B(n312), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U159 ( .A(n313), .B(n314), .Z(n312) );
  GTECH_XNOR2 U160 ( .A(n313), .B(n308), .Z(n311) );
  GTECH_AOI21 U161 ( .A(n315), .B(n316), .C(n317), .Z(n308) );
  GTECH_XOR2 U162 ( .A(n307), .B(n310), .Z(n313) );
  GTECH_NOT U163 ( .A(b[2]), .Z(n310) );
  GTECH_OAI21 U164 ( .A(n318), .B(n319), .C(n320), .Z(sum[1]) );
  GTECH_OAI21 U165 ( .A(n317), .B(n321), .C(n322), .Z(n320) );
  GTECH_OAI21 U166 ( .A(n323), .B(n324), .C(n325), .Z(n322) );
  GTECH_XNOR2 U167 ( .A(a[1]), .B(b[1]), .Z(n319) );
  GTECH_AOI21 U168 ( .A(n324), .B(n325), .C(n323), .Z(n318) );
  GTECH_NOT U169 ( .A(n316), .Z(n325) );
  GTECH_MUX2 U170 ( .A(n326), .B(n327), .S(n328), .Z(sum[15]) );
  GTECH_XOR2 U171 ( .A(n329), .B(n330), .Z(n327) );
  GTECH_AOI21 U172 ( .A(n331), .B(n332), .C(n333), .Z(n329) );
  GTECH_OA21 U173 ( .A(n332), .B(n331), .C(n334), .Z(n333) );
  GTECH_XOR2 U174 ( .A(n330), .B(n335), .Z(n326) );
  GTECH_XOR2 U175 ( .A(a[15]), .B(b[15]), .Z(n330) );
  GTECH_XNOR3 U176 ( .A(n334), .B(a[14]), .C(n336), .Z(sum[14]) );
  GTECH_OAI21 U177 ( .A(n337), .B(n328), .C(n332), .Z(n336) );
  GTECH_AOI21 U178 ( .A(n338), .B(n339), .C(n340), .Z(n332) );
  GTECH_NOT U179 ( .A(n341), .Z(n338) );
  GTECH_NOT U180 ( .A(b[14]), .Z(n334) );
  GTECH_MUX2 U181 ( .A(n342), .B(n343), .S(n328), .Z(sum[13]) );
  GTECH_XNOR2 U182 ( .A(n344), .B(n345), .Z(n343) );
  GTECH_NOT U183 ( .A(n339), .Z(n344) );
  GTECH_XOR2 U184 ( .A(n345), .B(n346), .Z(n342) );
  GTECH_NOT U185 ( .A(n347), .Z(n346) );
  GTECH_NOR2 U186 ( .A(n341), .B(n340), .Z(n345) );
  GTECH_NAND2 U187 ( .A(n348), .B(n349), .Z(sum[12]) );
  GTECH_OAI21 U188 ( .A(n339), .B(n347), .C(n350), .Z(n349) );
  GTECH_MUX2 U189 ( .A(n351), .B(n352), .S(n270), .Z(sum[11]) );
  GTECH_XNOR2 U190 ( .A(n353), .B(n354), .Z(n352) );
  GTECH_XOR2 U191 ( .A(n355), .B(n353), .Z(n351) );
  GTECH_XOR2 U192 ( .A(a[11]), .B(b[11]), .Z(n353) );
  GTECH_OA21 U193 ( .A(a[10]), .B(n356), .C(n357), .Z(n355) );
  GTECH_NOT U194 ( .A(n358), .Z(n357) );
  GTECH_AOI21 U195 ( .A(n356), .B(a[10]), .C(b[10]), .Z(n358) );
  GTECH_XNOR3 U196 ( .A(b[10]), .B(a[10]), .C(n359), .Z(sum[10]) );
  GTECH_AOI21 U197 ( .A(n360), .B(n270), .C(n356), .Z(n359) );
  GTECH_OAI21 U198 ( .A(n274), .B(n273), .C(n275), .Z(n356) );
  GTECH_NAND2 U199 ( .A(n361), .B(n362), .Z(sum[0]) );
  GTECH_OAI21 U200 ( .A(n316), .B(n323), .C(cin), .Z(n362) );
  GTECH_OAI21 U201 ( .A(n363), .B(n328), .C(n348), .Z(cout) );
  GTECH_OR3 U202 ( .A(n347), .B(n339), .C(n350), .Z(n348) );
  GTECH_NOT U203 ( .A(n328), .Z(n350) );
  GTECH_AND2 U204 ( .A(b[12]), .B(a[12]), .Z(n339) );
  GTECH_MUX2 U205 ( .A(n276), .B(n364), .S(n270), .Z(n328) );
  GTECH_MUX2 U206 ( .A(n365), .B(n301), .S(n279), .Z(n270) );
  GTECH_NOT U207 ( .A(n296), .Z(n279) );
  GTECH_OAI21 U208 ( .A(n366), .B(n324), .C(n361), .Z(n296) );
  GTECH_OR3 U209 ( .A(n323), .B(cin), .C(n316), .Z(n361) );
  GTECH_AND2 U210 ( .A(b[0]), .B(a[0]), .Z(n316) );
  GTECH_NOT U211 ( .A(cin), .Z(n324) );
  GTECH_AOI21 U212 ( .A(n305), .B(a[3]), .C(n367), .Z(n366) );
  GTECH_OA21 U213 ( .A(a[3]), .B(n305), .C(b[3]), .Z(n367) );
  GTECH_OAI21 U214 ( .A(n368), .B(n307), .C(n369), .Z(n305) );
  GTECH_OAI21 U215 ( .A(a[2]), .B(n314), .C(b[2]), .Z(n369) );
  GTECH_NOT U216 ( .A(n368), .Z(n314) );
  GTECH_NOT U217 ( .A(a[2]), .Z(n307) );
  GTECH_AOI21 U218 ( .A(n370), .B(n315), .C(n317), .Z(n368) );
  GTECH_AND2 U219 ( .A(b[1]), .B(a[1]), .Z(n317) );
  GTECH_NOT U220 ( .A(n321), .Z(n315) );
  GTECH_NOR2 U221 ( .A(a[1]), .B(b[1]), .Z(n321) );
  GTECH_NOT U222 ( .A(n323), .Z(n370) );
  GTECH_NOR2 U223 ( .A(a[0]), .B(b[0]), .Z(n323) );
  GTECH_XOR2 U224 ( .A(n298), .B(n299), .Z(n301) );
  GTECH_NOT U225 ( .A(b[4]), .Z(n299) );
  GTECH_AOI21 U226 ( .A(n371), .B(n286), .C(n372), .Z(n365) );
  GTECH_AOI21 U227 ( .A(n373), .B(a[7]), .C(b[7]), .Z(n372) );
  GTECH_NOT U228 ( .A(n286), .Z(n373) );
  GTECH_OA21 U229 ( .A(n288), .B(n282), .C(n374), .Z(n286) );
  GTECH_OAI21 U230 ( .A(a[6]), .B(n375), .C(b[6]), .Z(n374) );
  GTECH_NOT U231 ( .A(n288), .Z(n375) );
  GTECH_NOT U232 ( .A(a[6]), .Z(n282) );
  GTECH_AOI21 U233 ( .A(n297), .B(n289), .C(n291), .Z(n288) );
  GTECH_AND2 U234 ( .A(b[5]), .B(a[5]), .Z(n291) );
  GTECH_OR2 U235 ( .A(b[5]), .B(a[5]), .Z(n289) );
  GTECH_OR_NOT U236 ( .A(b[4]), .B(n298), .Z(n297) );
  GTECH_NOT U237 ( .A(a[4]), .Z(n298) );
  GTECH_NOT U238 ( .A(a[7]), .Z(n371) );
  GTECH_OAI21 U239 ( .A(a[11]), .B(n376), .C(n377), .Z(n364) );
  GTECH_NOT U240 ( .A(n378), .Z(n377) );
  GTECH_AOI21 U241 ( .A(n376), .B(a[11]), .C(b[11]), .Z(n378) );
  GTECH_NOT U242 ( .A(n354), .Z(n376) );
  GTECH_AOI21 U243 ( .A(n360), .B(a[10]), .C(n379), .Z(n354) );
  GTECH_OA21 U244 ( .A(a[10]), .B(n360), .C(b[10]), .Z(n379) );
  GTECH_OAI21 U245 ( .A(n272), .B(n274), .C(n275), .Z(n360) );
  GTECH_NAND2 U246 ( .A(b[9]), .B(a[9]), .Z(n275) );
  GTECH_NOR2 U247 ( .A(b[9]), .B(a[9]), .Z(n274) );
  GTECH_OR_NOT U248 ( .A(n272), .B(n273), .Z(n276) );
  GTECH_NAND2 U249 ( .A(b[8]), .B(a[8]), .Z(n273) );
  GTECH_NOR2 U250 ( .A(a[8]), .B(b[8]), .Z(n272) );
  GTECH_AOI21 U251 ( .A(n335), .B(a[15]), .C(n380), .Z(n363) );
  GTECH_OA21 U252 ( .A(a[15]), .B(n335), .C(b[15]), .Z(n380) );
  GTECH_OAI21 U253 ( .A(n337), .B(n331), .C(n381), .Z(n335) );
  GTECH_OAI21 U254 ( .A(a[14]), .B(n382), .C(b[14]), .Z(n381) );
  GTECH_NOT U255 ( .A(n337), .Z(n382) );
  GTECH_NOT U256 ( .A(a[14]), .Z(n331) );
  GTECH_OA21 U257 ( .A(n341), .B(n347), .C(n383), .Z(n337) );
  GTECH_NOT U258 ( .A(n340), .Z(n383) );
  GTECH_AND2 U259 ( .A(b[13]), .B(a[13]), .Z(n340) );
  GTECH_NOR2 U260 ( .A(b[12]), .B(a[12]), .Z(n347) );
  GTECH_NOR2 U261 ( .A(b[13]), .B(a[13]), .Z(n341) );
endmodule

