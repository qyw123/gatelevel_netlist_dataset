
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383;

  GTECH_MUX2 U138 ( .A(n277), .B(n278), .S(n279), .Z(sum[9]) );
  GTECH_OA21 U139 ( .A(n280), .B(n281), .C(n282), .Z(n279) );
  GTECH_OR_NOT U140 ( .A(n283), .B(n284), .Z(n278) );
  GTECH_XOR2 U141 ( .A(b[9]), .B(a[9]), .Z(n277) );
  GTECH_NAND2 U142 ( .A(n285), .B(n286), .Z(sum[8]) );
  GTECH_OAI21 U143 ( .A(n287), .B(n280), .C(n281), .Z(n285) );
  GTECH_MUX2 U144 ( .A(n288), .B(n289), .S(n290), .Z(sum[7]) );
  GTECH_XOR2 U145 ( .A(n291), .B(n292), .Z(n289) );
  GTECH_XNOR2 U146 ( .A(n291), .B(n293), .Z(n288) );
  GTECH_AND_NOT U147 ( .A(n294), .B(n295), .Z(n293) );
  GTECH_OAI21 U148 ( .A(b[6]), .B(a[6]), .C(n296), .Z(n294) );
  GTECH_XOR2 U149 ( .A(a[7]), .B(b[7]), .Z(n291) );
  GTECH_AO21 U150 ( .A(n297), .B(n295), .C(n298), .Z(sum[6]) );
  GTECH_NOT U151 ( .A(n299), .Z(n298) );
  GTECH_MUX2 U152 ( .A(n300), .B(n301), .S(b[6]), .Z(n299) );
  GTECH_OR_NOT U153 ( .A(n297), .B(n302), .Z(n301) );
  GTECH_XOR2 U154 ( .A(n302), .B(n297), .Z(n300) );
  GTECH_NOT U155 ( .A(a[6]), .Z(n302) );
  GTECH_AO21 U156 ( .A(n290), .B(n303), .C(n296), .Z(n297) );
  GTECH_AOI21 U157 ( .A(n304), .B(n305), .C(n306), .Z(n296) );
  GTECH_MUX2 U158 ( .A(n307), .B(n308), .S(n309), .Z(sum[5]) );
  GTECH_AND_NOT U159 ( .A(n305), .B(n306), .Z(n309) );
  GTECH_OAI21 U160 ( .A(n310), .B(n290), .C(n311), .Z(n308) );
  GTECH_AO21 U161 ( .A(n311), .B(n290), .C(n310), .Z(n307) );
  GTECH_NOT U162 ( .A(n304), .Z(n310) );
  GTECH_XOR2 U163 ( .A(n312), .B(n290), .Z(sum[4]) );
  GTECH_MUX2 U164 ( .A(n313), .B(n314), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U165 ( .A(n315), .B(n316), .Z(n314) );
  GTECH_XOR2 U166 ( .A(n317), .B(n315), .Z(n313) );
  GTECH_XOR2 U167 ( .A(a[3]), .B(b[3]), .Z(n315) );
  GTECH_ADD_ABC U168 ( .A(a[2]), .B(n318), .C(b[2]), .COUT(n317) );
  GTECH_MUX2 U169 ( .A(n319), .B(n320), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U170 ( .A(n321), .B(n322), .Z(n320) );
  GTECH_XOR2 U171 ( .A(n318), .B(n322), .Z(n319) );
  GTECH_XOR2 U172 ( .A(a[2]), .B(b[2]), .Z(n322) );
  GTECH_OA21 U173 ( .A(n323), .B(n324), .C(n325), .Z(n318) );
  GTECH_MUX2 U174 ( .A(n326), .B(n327), .S(n328), .Z(sum[1]) );
  GTECH_AND_NOT U175 ( .A(n325), .B(n323), .Z(n328) );
  GTECH_OAI21 U176 ( .A(cin), .B(n324), .C(n329), .Z(n327) );
  GTECH_AO21 U177 ( .A(n329), .B(cin), .C(n324), .Z(n326) );
  GTECH_MUX2 U178 ( .A(n330), .B(n331), .S(n332), .Z(sum[15]) );
  GTECH_XOR2 U179 ( .A(n333), .B(n334), .Z(n331) );
  GTECH_OA21 U180 ( .A(n335), .B(n336), .C(n337), .Z(n334) );
  GTECH_XNOR2 U181 ( .A(n333), .B(n338), .Z(n330) );
  GTECH_XNOR2 U182 ( .A(a[15]), .B(b[15]), .Z(n333) );
  GTECH_MUX2 U183 ( .A(n339), .B(n340), .S(n341), .Z(sum[14]) );
  GTECH_OA21 U184 ( .A(n332), .B(n342), .C(n336), .Z(n341) );
  GTECH_OAI21 U185 ( .A(n343), .B(n344), .C(n345), .Z(n336) );
  GTECH_XOR2 U186 ( .A(b[14]), .B(a[14]), .Z(n340) );
  GTECH_OR_NOT U187 ( .A(n335), .B(n337), .Z(n339) );
  GTECH_MUX2 U188 ( .A(n346), .B(n347), .S(n348), .Z(sum[13]) );
  GTECH_MUX2 U189 ( .A(n349), .B(n350), .S(n351), .Z(n347) );
  GTECH_MUX2 U190 ( .A(n350), .B(n349), .S(n343), .Z(n346) );
  GTECH_OR_NOT U191 ( .A(n344), .B(n345), .Z(n349) );
  GTECH_XOR2 U192 ( .A(a[13]), .B(b[13]), .Z(n350) );
  GTECH_XOR2 U193 ( .A(n352), .B(n348), .Z(sum[12]) );
  GTECH_NOT U194 ( .A(n332), .Z(n348) );
  GTECH_MUX2 U195 ( .A(n353), .B(n354), .S(n355), .Z(sum[11]) );
  GTECH_XNOR2 U196 ( .A(n356), .B(n357), .Z(n354) );
  GTECH_OA21 U197 ( .A(n358), .B(n359), .C(n360), .Z(n357) );
  GTECH_XOR2 U198 ( .A(n356), .B(n361), .Z(n353) );
  GTECH_XOR2 U199 ( .A(a[11]), .B(b[11]), .Z(n356) );
  GTECH_MUX2 U200 ( .A(n362), .B(n363), .S(n364), .Z(sum[10]) );
  GTECH_OA21 U201 ( .A(n355), .B(n365), .C(n359), .Z(n364) );
  GTECH_OAI21 U202 ( .A(n283), .B(n280), .C(n284), .Z(n359) );
  GTECH_XOR2 U203 ( .A(b[10]), .B(a[10]), .Z(n363) );
  GTECH_OR_NOT U204 ( .A(n358), .B(n360), .Z(n362) );
  GTECH_XNOR2 U205 ( .A(n366), .B(n367), .Z(sum[0]) );
  GTECH_MUX2 U206 ( .A(n368), .B(n352), .S(n332), .Z(cout) );
  GTECH_OA21 U207 ( .A(n369), .B(n355), .C(n286), .Z(n332) );
  GTECH_OR3 U208 ( .A(n280), .B(n287), .C(n281), .Z(n286) );
  GTECH_AND2 U209 ( .A(b[8]), .B(a[8]), .Z(n280) );
  GTECH_NOT U210 ( .A(n281), .Z(n355) );
  GTECH_MUX2 U211 ( .A(n312), .B(n370), .S(n290), .Z(n281) );
  GTECH_MUX2 U212 ( .A(n371), .B(n367), .S(n366), .Z(n290) );
  GTECH_NOT U213 ( .A(cin), .Z(n366) );
  GTECH_AND_NOT U214 ( .A(n329), .B(n324), .Z(n367) );
  GTECH_AND2 U215 ( .A(b[0]), .B(a[0]), .Z(n324) );
  GTECH_AO21 U216 ( .A(n316), .B(a[3]), .C(n372), .Z(n371) );
  GTECH_OA21 U217 ( .A(a[3]), .B(n316), .C(b[3]), .Z(n372) );
  GTECH_ADD_ABC U218 ( .A(n321), .B(a[2]), .C(b[2]), .COUT(n316) );
  GTECH_OA21 U219 ( .A(n323), .B(n329), .C(n325), .Z(n321) );
  GTECH_OR_NOT U220 ( .A(a[1]), .B(n373), .Z(n325) );
  GTECH_NOT U221 ( .A(b[1]), .Z(n373) );
  GTECH_NOT U222 ( .A(n374), .Z(n329) );
  GTECH_NOR2 U223 ( .A(b[0]), .B(a[0]), .Z(n374) );
  GTECH_AND2 U224 ( .A(a[1]), .B(b[1]), .Z(n323) );
  GTECH_OA21 U225 ( .A(a[7]), .B(n292), .C(n375), .Z(n370) );
  GTECH_AO21 U226 ( .A(n292), .B(a[7]), .C(b[7]), .Z(n375) );
  GTECH_OR_NOT U227 ( .A(n295), .B(n376), .Z(n292) );
  GTECH_OAI21 U228 ( .A(a[6]), .B(b[6]), .C(n303), .Z(n376) );
  GTECH_AOI21 U229 ( .A(n305), .B(n377), .C(n306), .Z(n303) );
  GTECH_NOR2 U230 ( .A(b[5]), .B(a[5]), .Z(n306) );
  GTECH_NAND2 U231 ( .A(b[5]), .B(a[5]), .Z(n305) );
  GTECH_AND2 U232 ( .A(b[6]), .B(a[6]), .Z(n295) );
  GTECH_AND2 U233 ( .A(n311), .B(n304), .Z(n312) );
  GTECH_NAND2 U234 ( .A(b[4]), .B(a[4]), .Z(n304) );
  GTECH_NOT U235 ( .A(n377), .Z(n311) );
  GTECH_NOR2 U236 ( .A(b[4]), .B(a[4]), .Z(n377) );
  GTECH_AOI21 U237 ( .A(n361), .B(a[11]), .C(n378), .Z(n369) );
  GTECH_OA21 U238 ( .A(a[11]), .B(n361), .C(b[11]), .Z(n378) );
  GTECH_OAI21 U239 ( .A(n358), .B(n365), .C(n360), .Z(n361) );
  GTECH_NAND2 U240 ( .A(a[10]), .B(b[10]), .Z(n360) );
  GTECH_OAI21 U241 ( .A(n283), .B(n282), .C(n284), .Z(n365) );
  GTECH_OR_NOT U242 ( .A(b[9]), .B(n379), .Z(n284) );
  GTECH_NOT U243 ( .A(a[9]), .Z(n379) );
  GTECH_NOT U244 ( .A(n287), .Z(n282) );
  GTECH_NOR2 U245 ( .A(b[8]), .B(a[8]), .Z(n287) );
  GTECH_AND2 U246 ( .A(b[9]), .B(a[9]), .Z(n283) );
  GTECH_NOR2 U247 ( .A(b[10]), .B(a[10]), .Z(n358) );
  GTECH_AND_NOT U248 ( .A(n380), .B(n343), .Z(n352) );
  GTECH_AND2 U249 ( .A(b[12]), .B(a[12]), .Z(n343) );
  GTECH_AO21 U250 ( .A(n338), .B(a[15]), .C(n381), .Z(n368) );
  GTECH_OA21 U251 ( .A(a[15]), .B(n338), .C(b[15]), .Z(n381) );
  GTECH_OAI21 U252 ( .A(n335), .B(n342), .C(n337), .Z(n338) );
  GTECH_OR_NOT U253 ( .A(n382), .B(b[14]), .Z(n337) );
  GTECH_NOT U254 ( .A(a[14]), .Z(n382) );
  GTECH_OAI21 U255 ( .A(n344), .B(n380), .C(n345), .Z(n342) );
  GTECH_OR_NOT U256 ( .A(a[13]), .B(n383), .Z(n345) );
  GTECH_NOT U257 ( .A(n351), .Z(n380) );
  GTECH_NOR2 U258 ( .A(b[12]), .B(a[12]), .Z(n351) );
  GTECH_AND_NOT U259 ( .A(a[13]), .B(n383), .Z(n344) );
  GTECH_NOT U260 ( .A(b[13]), .Z(n383) );
  GTECH_NOR2 U261 ( .A(a[14]), .B(b[14]), .Z(n335) );
endmodule

