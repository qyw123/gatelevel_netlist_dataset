
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128;

  GTECH_XOR2 U81 ( .A(n62), .B(n63), .Z(sum[9]) );
  GTECH_XNOR2 U82 ( .A(n64), .B(n65), .Z(sum[8]) );
  GTECH_XOR2 U83 ( .A(n66), .B(n67), .Z(sum[7]) );
  GTECH_OA21 U84 ( .A(n68), .B(n69), .C(n70), .Z(n67) );
  GTECH_XOR2 U85 ( .A(n69), .B(n68), .Z(sum[6]) );
  GTECH_OA21 U86 ( .A(n71), .B(n72), .C(n73), .Z(n68) );
  GTECH_XOR2 U87 ( .A(n72), .B(n71), .Z(sum[5]) );
  GTECH_OA21 U88 ( .A(n74), .B(n75), .C(n76), .Z(n71) );
  GTECH_XOR2 U89 ( .A(n75), .B(n74), .Z(sum[4]) );
  GTECH_XOR2 U90 ( .A(n77), .B(n78), .Z(sum[3]) );
  GTECH_OA21 U91 ( .A(n79), .B(n80), .C(n81), .Z(n78) );
  GTECH_XOR2 U92 ( .A(n80), .B(n79), .Z(sum[2]) );
  GTECH_OA21 U93 ( .A(n82), .B(n83), .C(n84), .Z(n79) );
  GTECH_XOR2 U94 ( .A(n83), .B(n82), .Z(sum[1]) );
  GTECH_OA21 U95 ( .A(n85), .B(n86), .C(n87), .Z(n82) );
  GTECH_XOR2 U96 ( .A(n88), .B(n89), .Z(sum[15]) );
  GTECH_OA21 U97 ( .A(n90), .B(n91), .C(n92), .Z(n89) );
  GTECH_XOR2 U98 ( .A(n91), .B(n90), .Z(sum[14]) );
  GTECH_OA21 U99 ( .A(n93), .B(n94), .C(n95), .Z(n90) );
  GTECH_XOR2 U100 ( .A(n94), .B(n93), .Z(sum[13]) );
  GTECH_OA21 U101 ( .A(n96), .B(n97), .C(n98), .Z(n93) );
  GTECH_XNOR2 U102 ( .A(cout), .B(n97), .Z(sum[12]) );
  GTECH_XNOR2 U103 ( .A(n99), .B(n100), .Z(sum[11]) );
  GTECH_OAI21 U104 ( .A(n101), .B(n102), .C(n103), .Z(n99) );
  GTECH_XOR2 U105 ( .A(n102), .B(n101), .Z(sum[10]) );
  GTECH_AOI21 U106 ( .A(n63), .B(n62), .C(n104), .Z(n101) );
  GTECH_OAI21 U107 ( .A(n65), .B(n105), .C(n106), .Z(n63) );
  GTECH_NOT U108 ( .A(n64), .Z(n105) );
  GTECH_XNOR2 U109 ( .A(cin), .B(n85), .Z(sum[0]) );
  GTECH_NOT U110 ( .A(n96), .Z(cout) );
  GTECH_OA21 U111 ( .A(n65), .B(n107), .C(n108), .Z(n96) );
  GTECH_OA21 U112 ( .A(n74), .B(n109), .C(n110), .Z(n65) );
  GTECH_OA21 U113 ( .A(n111), .B(n86), .C(n112), .Z(n74) );
  GTECH_NOT U114 ( .A(cin), .Z(n86) );
  GTECH_NOR3 U115 ( .A(n109), .B(n111), .C(n107), .Z(Pm) );
  GTECH_OR5 U116 ( .A(n77), .B(n83), .C(n80), .D(n85), .E(n113), .Z(n111) );
  GTECH_OAI21 U117 ( .A(b[0]), .B(a[0]), .C(n87), .Z(n85) );
  GTECH_OAI21 U118 ( .A(n114), .B(n107), .C(n108), .Z(Gm) );
  GTECH_AOI2N2 U119 ( .A(b[15]), .B(a[15]), .C(n115), .D(n88), .Z(n108) );
  GTECH_OA21 U120 ( .A(n116), .B(n91), .C(n92), .Z(n115) );
  GTECH_OA21 U121 ( .A(n94), .B(n98), .C(n95), .Z(n116) );
  GTECH_NAND2 U122 ( .A(b[13]), .B(a[13]), .Z(n95) );
  GTECH_OR4 U123 ( .A(n97), .B(n91), .C(n88), .D(n94), .Z(n107) );
  GTECH_XNOR2 U124 ( .A(a[13]), .B(b[13]), .Z(n94) );
  GTECH_XNOR2 U125 ( .A(a[15]), .B(b[15]), .Z(n88) );
  GTECH_OAI21 U126 ( .A(b[14]), .B(a[14]), .C(n92), .Z(n91) );
  GTECH_NAND2 U127 ( .A(b[14]), .B(a[14]), .Z(n92) );
  GTECH_OAI21 U128 ( .A(b[12]), .B(a[12]), .C(n98), .Z(n97) );
  GTECH_NAND2 U129 ( .A(a[12]), .B(b[12]), .Z(n98) );
  GTECH_OA21 U130 ( .A(n112), .B(n109), .C(n110), .Z(n114) );
  GTECH_OA21 U131 ( .A(n117), .B(n100), .C(n118), .Z(n110) );
  GTECH_OA21 U132 ( .A(n119), .B(n102), .C(n103), .Z(n117) );
  GTECH_NOT U133 ( .A(n120), .Z(n102) );
  GTECH_AOI21 U134 ( .A(n62), .B(n121), .C(n104), .Z(n119) );
  GTECH_AND2 U135 ( .A(a[9]), .B(b[9]), .Z(n104) );
  GTECH_NAND4 U136 ( .A(n64), .B(n122), .C(n120), .D(n62), .Z(n109) );
  GTECH_XOR2 U137 ( .A(a[9]), .B(b[9]), .Z(n62) );
  GTECH_OA21 U138 ( .A(b[10]), .B(a[10]), .C(n103), .Z(n120) );
  GTECH_NAND2 U139 ( .A(b[10]), .B(a[10]), .Z(n103) );
  GTECH_NOT U140 ( .A(n100), .Z(n122) );
  GTECH_OAI21 U141 ( .A(b[11]), .B(a[11]), .C(n118), .Z(n100) );
  GTECH_NAND2 U142 ( .A(a[11]), .B(b[11]), .Z(n118) );
  GTECH_OA21 U143 ( .A(b[8]), .B(a[8]), .C(n106), .Z(n64) );
  GTECH_NOT U144 ( .A(n121), .Z(n106) );
  GTECH_AND2 U145 ( .A(a[8]), .B(b[8]), .Z(n121) );
  GTECH_AOI21 U146 ( .A(b[7]), .B(a[7]), .C(n123), .Z(n112) );
  GTECH_OAI22 U147 ( .A(n124), .B(n113), .C(n125), .D(n66), .Z(n123) );
  GTECH_OA21 U148 ( .A(n126), .B(n69), .C(n70), .Z(n125) );
  GTECH_OA21 U149 ( .A(n72), .B(n76), .C(n73), .Z(n126) );
  GTECH_OR4 U150 ( .A(n75), .B(n69), .C(n72), .D(n66), .Z(n113) );
  GTECH_XNOR2 U151 ( .A(a[7]), .B(b[7]), .Z(n66) );
  GTECH_OAI21 U152 ( .A(b[5]), .B(a[5]), .C(n73), .Z(n72) );
  GTECH_NAND2 U153 ( .A(b[5]), .B(a[5]), .Z(n73) );
  GTECH_OAI21 U154 ( .A(b[6]), .B(a[6]), .C(n70), .Z(n69) );
  GTECH_NAND2 U155 ( .A(b[6]), .B(a[6]), .Z(n70) );
  GTECH_OAI21 U156 ( .A(b[4]), .B(a[4]), .C(n76), .Z(n75) );
  GTECH_NAND2 U157 ( .A(b[4]), .B(a[4]), .Z(n76) );
  GTECH_AOI2N2 U158 ( .A(b[3]), .B(a[3]), .C(n127), .D(n77), .Z(n124) );
  GTECH_XNOR2 U159 ( .A(a[3]), .B(b[3]), .Z(n77) );
  GTECH_OA21 U160 ( .A(n128), .B(n80), .C(n81), .Z(n127) );
  GTECH_OAI21 U161 ( .A(b[2]), .B(a[2]), .C(n81), .Z(n80) );
  GTECH_NAND2 U162 ( .A(b[2]), .B(a[2]), .Z(n81) );
  GTECH_OA21 U163 ( .A(n83), .B(n87), .C(n84), .Z(n128) );
  GTECH_NAND2 U164 ( .A(a[1]), .B(b[1]), .Z(n84) );
  GTECH_NAND2 U165 ( .A(a[0]), .B(b[0]), .Z(n87) );
  GTECH_XNOR2 U166 ( .A(a[1]), .B(b[1]), .Z(n83) );
endmodule

