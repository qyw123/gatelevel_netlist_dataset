
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391;

  GTECH_MUX2 U149 ( .A(n288), .B(n289), .S(n290), .Z(sum[9]) );
  GTECH_XOR2 U150 ( .A(n291), .B(n292), .Z(n289) );
  GTECH_XNOR2 U151 ( .A(n293), .B(n291), .Z(n288) );
  GTECH_NOR2 U152 ( .A(n294), .B(n295), .Z(n291) );
  GTECH_XNOR2 U153 ( .A(n296), .B(n297), .Z(sum[8]) );
  GTECH_MUX2 U154 ( .A(n298), .B(n299), .S(n300), .Z(sum[7]) );
  GTECH_XOR2 U155 ( .A(n301), .B(n302), .Z(n299) );
  GTECH_OA21 U156 ( .A(n303), .B(n304), .C(n305), .Z(n302) );
  GTECH_XNOR2 U157 ( .A(n301), .B(n306), .Z(n298) );
  GTECH_XNOR2 U158 ( .A(a[7]), .B(b[7]), .Z(n301) );
  GTECH_MUX2 U159 ( .A(n307), .B(n308), .S(n309), .Z(sum[6]) );
  GTECH_OA21 U160 ( .A(n310), .B(n300), .C(n304), .Z(n309) );
  GTECH_AOI2N2 U161 ( .A(a[5]), .B(b[5]), .C(n311), .D(n312), .Z(n304) );
  GTECH_XOR2 U162 ( .A(b[6]), .B(a[6]), .Z(n308) );
  GTECH_NOT U163 ( .A(n313), .Z(n307) );
  GTECH_AND_NOT U164 ( .A(n305), .B(n303), .Z(n313) );
  GTECH_MUX2 U165 ( .A(n314), .B(n315), .S(n316), .Z(sum[5]) );
  GTECH_AOI21 U166 ( .A(a[5]), .B(b[5]), .C(n311), .Z(n316) );
  GTECH_OAI21 U167 ( .A(n317), .B(n318), .C(n319), .Z(n315) );
  GTECH_OAI21 U168 ( .A(n320), .B(n300), .C(n312), .Z(n314) );
  GTECH_XOR2 U169 ( .A(n300), .B(n321), .Z(sum[4]) );
  GTECH_MUX2 U170 ( .A(n322), .B(n323), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U171 ( .A(n324), .B(n325), .Z(n323) );
  GTECH_XOR2 U172 ( .A(n324), .B(n326), .Z(n322) );
  GTECH_AND2 U173 ( .A(n327), .B(n328), .Z(n326) );
  GTECH_OAI21 U174 ( .A(b[2]), .B(a[2]), .C(n329), .Z(n327) );
  GTECH_XNOR2 U175 ( .A(a[3]), .B(b[3]), .Z(n324) );
  GTECH_MUX2 U176 ( .A(n330), .B(n331), .S(n332), .Z(sum[2]) );
  GTECH_MUX2 U177 ( .A(n333), .B(n334), .S(n329), .Z(n331) );
  GTECH_OAI21 U178 ( .A(n335), .B(n336), .C(n337), .Z(n329) );
  GTECH_MUX2 U179 ( .A(n333), .B(n334), .S(n338), .Z(n330) );
  GTECH_OAI21 U180 ( .A(b[2]), .B(a[2]), .C(n328), .Z(n334) );
  GTECH_XOR2 U181 ( .A(a[2]), .B(b[2]), .Z(n333) );
  GTECH_MUX2 U182 ( .A(n339), .B(n340), .S(n341), .Z(sum[1]) );
  GTECH_AND_NOT U183 ( .A(n337), .B(n335), .Z(n341) );
  GTECH_AO21 U184 ( .A(n332), .B(n336), .C(n342), .Z(n340) );
  GTECH_OAI21 U185 ( .A(n342), .B(n332), .C(n336), .Z(n339) );
  GTECH_NAND2 U186 ( .A(a[0]), .B(b[0]), .Z(n336) );
  GTECH_MUX2 U187 ( .A(n343), .B(n344), .S(n345), .Z(sum[15]) );
  GTECH_XOR2 U188 ( .A(n346), .B(n347), .Z(n344) );
  GTECH_OA21 U189 ( .A(n348), .B(n349), .C(n350), .Z(n347) );
  GTECH_XNOR2 U190 ( .A(n346), .B(n351), .Z(n343) );
  GTECH_XNOR2 U191 ( .A(a[15]), .B(b[15]), .Z(n346) );
  GTECH_MUX2 U192 ( .A(n352), .B(n353), .S(n354), .Z(sum[14]) );
  GTECH_OA21 U193 ( .A(n355), .B(n345), .C(n349), .Z(n354) );
  GTECH_AOI2N2 U194 ( .A(a[13]), .B(b[13]), .C(n356), .D(n357), .Z(n349) );
  GTECH_XOR2 U195 ( .A(b[14]), .B(a[14]), .Z(n353) );
  GTECH_NOT U196 ( .A(n358), .Z(n352) );
  GTECH_AND_NOT U197 ( .A(n350), .B(n348), .Z(n358) );
  GTECH_MUX2 U198 ( .A(n359), .B(n360), .S(n345), .Z(sum[13]) );
  GTECH_XNOR2 U199 ( .A(n361), .B(n357), .Z(n360) );
  GTECH_XOR2 U200 ( .A(n361), .B(n362), .Z(n359) );
  GTECH_AOI21 U201 ( .A(a[13]), .B(b[13]), .C(n356), .Z(n361) );
  GTECH_NAND2 U202 ( .A(n363), .B(n364), .Z(sum[12]) );
  GTECH_AO21 U203 ( .A(n357), .B(n362), .C(n345), .Z(n363) );
  GTECH_MUX2 U204 ( .A(n365), .B(n366), .S(n297), .Z(sum[11]) );
  GTECH_XOR2 U205 ( .A(n367), .B(n368), .Z(n366) );
  GTECH_OA21 U206 ( .A(n369), .B(n370), .C(n371), .Z(n368) );
  GTECH_XNOR2 U207 ( .A(n367), .B(n372), .Z(n365) );
  GTECH_XNOR2 U208 ( .A(a[11]), .B(b[11]), .Z(n367) );
  GTECH_MUX2 U209 ( .A(n373), .B(n374), .S(n297), .Z(sum[10]) );
  GTECH_XNOR2 U210 ( .A(n370), .B(n375), .Z(n374) );
  GTECH_AOI21 U211 ( .A(n376), .B(n377), .C(n295), .Z(n370) );
  GTECH_XNOR2 U212 ( .A(n375), .B(n378), .Z(n373) );
  GTECH_AND_NOT U213 ( .A(n371), .B(n369), .Z(n375) );
  GTECH_XNOR2 U214 ( .A(n332), .B(n379), .Z(sum[0]) );
  GTECH_NOT U215 ( .A(cin), .Z(n332) );
  GTECH_OAI21 U216 ( .A(n380), .B(n345), .C(n364), .Z(cout) );
  GTECH_NAND3 U217 ( .A(n357), .B(n362), .C(n345), .Z(n364) );
  GTECH_NOT U218 ( .A(n381), .Z(n362) );
  GTECH_NAND2 U219 ( .A(a[12]), .B(b[12]), .Z(n357) );
  GTECH_NOT U220 ( .A(n382), .Z(n345) );
  GTECH_MUX2 U221 ( .A(n296), .B(n383), .S(n290), .Z(n382) );
  GTECH_NOT U222 ( .A(n297), .Z(n290) );
  GTECH_MUX2 U223 ( .A(n384), .B(n321), .S(n300), .Z(n297) );
  GTECH_NOT U224 ( .A(n318), .Z(n300) );
  GTECH_MUX2 U225 ( .A(n379), .B(n385), .S(cin), .Z(n318) );
  GTECH_OA21 U226 ( .A(a[3]), .B(n325), .C(n386), .Z(n385) );
  GTECH_AO21 U227 ( .A(n325), .B(a[3]), .C(b[3]), .Z(n386) );
  GTECH_NAND2 U228 ( .A(n387), .B(n328), .Z(n325) );
  GTECH_NAND2 U229 ( .A(b[2]), .B(a[2]), .Z(n328) );
  GTECH_OAI21 U230 ( .A(a[2]), .B(b[2]), .C(n338), .Z(n387) );
  GTECH_OAI21 U231 ( .A(n342), .B(n335), .C(n337), .Z(n338) );
  GTECH_NAND2 U232 ( .A(b[1]), .B(a[1]), .Z(n337) );
  GTECH_NOR2 U233 ( .A(b[1]), .B(a[1]), .Z(n335) );
  GTECH_NOR2 U234 ( .A(b[0]), .B(a[0]), .Z(n342) );
  GTECH_XOR2 U235 ( .A(a[0]), .B(b[0]), .Z(n379) );
  GTECH_NAND2 U236 ( .A(n319), .B(n312), .Z(n321) );
  GTECH_NOT U237 ( .A(n317), .Z(n312) );
  GTECH_AND2 U238 ( .A(b[4]), .B(a[4]), .Z(n317) );
  GTECH_NOT U239 ( .A(n320), .Z(n319) );
  GTECH_AOI21 U240 ( .A(n306), .B(a[7]), .C(n388), .Z(n384) );
  GTECH_OA21 U241 ( .A(a[7]), .B(n306), .C(b[7]), .Z(n388) );
  GTECH_OAI21 U242 ( .A(n303), .B(n310), .C(n305), .Z(n306) );
  GTECH_NAND2 U243 ( .A(a[6]), .B(b[6]), .Z(n305) );
  GTECH_AOI2N2 U244 ( .A(a[5]), .B(b[5]), .C(n311), .D(n320), .Z(n310) );
  GTECH_NOR2 U245 ( .A(b[4]), .B(a[4]), .Z(n320) );
  GTECH_NOR2 U246 ( .A(a[5]), .B(b[5]), .Z(n311) );
  GTECH_NOR2 U247 ( .A(b[6]), .B(a[6]), .Z(n303) );
  GTECH_OA21 U248 ( .A(a[11]), .B(n372), .C(n389), .Z(n383) );
  GTECH_AO21 U249 ( .A(n372), .B(a[11]), .C(b[11]), .Z(n389) );
  GTECH_OAI21 U250 ( .A(n378), .B(n369), .C(n371), .Z(n372) );
  GTECH_NAND2 U251 ( .A(a[10]), .B(b[10]), .Z(n371) );
  GTECH_NOR2 U252 ( .A(a[10]), .B(b[10]), .Z(n369) );
  GTECH_AOI21 U253 ( .A(n376), .B(n292), .C(n295), .Z(n378) );
  GTECH_AND2 U254 ( .A(b[9]), .B(a[9]), .Z(n295) );
  GTECH_NOT U255 ( .A(n390), .Z(n292) );
  GTECH_NOT U256 ( .A(n294), .Z(n376) );
  GTECH_NOR2 U257 ( .A(a[9]), .B(b[9]), .Z(n294) );
  GTECH_AND_NOT U258 ( .A(n293), .B(n390), .Z(n296) );
  GTECH_NOR2 U259 ( .A(b[8]), .B(a[8]), .Z(n390) );
  GTECH_NOT U260 ( .A(n377), .Z(n293) );
  GTECH_AND2 U261 ( .A(b[8]), .B(a[8]), .Z(n377) );
  GTECH_AOI21 U262 ( .A(n351), .B(a[15]), .C(n391), .Z(n380) );
  GTECH_OA21 U263 ( .A(a[15]), .B(n351), .C(b[15]), .Z(n391) );
  GTECH_OAI21 U264 ( .A(n348), .B(n355), .C(n350), .Z(n351) );
  GTECH_NAND2 U265 ( .A(a[14]), .B(b[14]), .Z(n350) );
  GTECH_AOI2N2 U266 ( .A(a[13]), .B(b[13]), .C(n356), .D(n381), .Z(n355) );
  GTECH_NOR2 U267 ( .A(b[12]), .B(a[12]), .Z(n381) );
  GTECH_NOR2 U268 ( .A(a[13]), .B(b[13]), .Z(n356) );
  GTECH_NOR2 U269 ( .A(b[14]), .B(a[14]), .Z(n348) );
endmodule

