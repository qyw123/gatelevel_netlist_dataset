
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133;

  GTECH_XOR2 U87 ( .A(n68), .B(n69), .Z(sum[9]) );
  GTECH_XOR2 U88 ( .A(n70), .B(n71), .Z(sum[8]) );
  GTECH_XNOR2 U89 ( .A(n72), .B(n73), .Z(sum[7]) );
  GTECH_AOI21 U90 ( .A(n74), .B(n75), .C(n76), .Z(n73) );
  GTECH_XOR2 U91 ( .A(n74), .B(n75), .Z(sum[6]) );
  GTECH_AO22 U92 ( .A(b[5]), .B(a[5]), .C(n77), .D(n78), .Z(n74) );
  GTECH_XOR2 U93 ( .A(n78), .B(n77), .Z(sum[5]) );
  GTECH_AO22 U94 ( .A(a[4]), .B(b[4]), .C(n79), .D(n80), .Z(n77) );
  GTECH_XOR2 U95 ( .A(n80), .B(n79), .Z(sum[4]) );
  GTECH_NOT U96 ( .A(n81), .Z(n79) );
  GTECH_XNOR2 U97 ( .A(n82), .B(n83), .Z(sum[3]) );
  GTECH_AOI21 U98 ( .A(n84), .B(n85), .C(n86), .Z(n83) );
  GTECH_XOR2 U99 ( .A(n85), .B(n84), .Z(sum[2]) );
  GTECH_AO22 U100 ( .A(b[1]), .B(a[1]), .C(n87), .D(n88), .Z(n84) );
  GTECH_XOR2 U101 ( .A(n88), .B(n87), .Z(sum[1]) );
  GTECH_AO22 U102 ( .A(a[0]), .B(b[0]), .C(n89), .D(cin), .Z(n87) );
  GTECH_XNOR2 U103 ( .A(n90), .B(n91), .Z(sum[15]) );
  GTECH_OA21 U104 ( .A(n92), .B(n93), .C(n94), .Z(n91) );
  GTECH_XNOR2 U105 ( .A(n95), .B(n92), .Z(sum[14]) );
  GTECH_OA21 U106 ( .A(n96), .B(n97), .C(n98), .Z(n92) );
  GTECH_XOR2 U107 ( .A(n97), .B(n96), .Z(sum[13]) );
  GTECH_AOI21 U108 ( .A(cout), .B(n99), .C(n100), .Z(n96) );
  GTECH_NOT U109 ( .A(n101), .Z(n100) );
  GTECH_XOR2 U110 ( .A(cout), .B(n99), .Z(sum[12]) );
  GTECH_XOR2 U111 ( .A(n102), .B(n103), .Z(sum[11]) );
  GTECH_AO21 U112 ( .A(n104), .B(n105), .C(n106), .Z(n102) );
  GTECH_XOR2 U113 ( .A(n104), .B(n105), .Z(sum[10]) );
  GTECH_AO22 U114 ( .A(b[9]), .B(a[9]), .C(n69), .D(n68), .Z(n104) );
  GTECH_AO22 U115 ( .A(a[8]), .B(b[8]), .C(n71), .D(n70), .Z(n69) );
  GTECH_XNOR2 U116 ( .A(n107), .B(n89), .Z(sum[0]) );
  GTECH_OAI21 U117 ( .A(n108), .B(n109), .C(n110), .Z(cout) );
  GTECH_NOT U118 ( .A(n71), .Z(n108) );
  GTECH_OAI21 U119 ( .A(n81), .B(n111), .C(n112), .Z(n71) );
  GTECH_OA21 U120 ( .A(n113), .B(n107), .C(n114), .Z(n81) );
  GTECH_NOT U121 ( .A(cin), .Z(n107) );
  GTECH_NOR3 U122 ( .A(n111), .B(n113), .C(n109), .Z(Pm) );
  GTECH_NAND5 U123 ( .A(n85), .B(n88), .C(n82), .D(n115), .E(n89), .Z(n113) );
  GTECH_XOR2 U124 ( .A(a[0]), .B(b[0]), .Z(n89) );
  GTECH_OAI21 U125 ( .A(n116), .B(n109), .C(n110), .Z(Gm) );
  GTECH_AOI22 U126 ( .A(b[15]), .B(a[15]), .C(n117), .D(n90), .Z(n110) );
  GTECH_OAI21 U127 ( .A(n118), .B(n93), .C(n94), .Z(n117) );
  GTECH_OA21 U128 ( .A(n97), .B(n101), .C(n98), .Z(n118) );
  GTECH_NAND2 U129 ( .A(b[13]), .B(a[13]), .Z(n98) );
  GTECH_NOT U130 ( .A(n119), .Z(n97) );
  GTECH_NAND4 U131 ( .A(n99), .B(n95), .C(n90), .D(n119), .Z(n109) );
  GTECH_XOR2 U132 ( .A(a[13]), .B(b[13]), .Z(n119) );
  GTECH_XOR2 U133 ( .A(a[15]), .B(b[15]), .Z(n90) );
  GTECH_NOT U134 ( .A(n93), .Z(n95) );
  GTECH_OAI21 U135 ( .A(b[14]), .B(a[14]), .C(n94), .Z(n93) );
  GTECH_NAND2 U136 ( .A(b[14]), .B(a[14]), .Z(n94) );
  GTECH_OA21 U137 ( .A(b[12]), .B(a[12]), .C(n101), .Z(n99) );
  GTECH_NAND2 U138 ( .A(a[12]), .B(b[12]), .Z(n101) );
  GTECH_OA21 U139 ( .A(n114), .B(n111), .C(n112), .Z(n116) );
  GTECH_AOI21 U140 ( .A(n120), .B(n103), .C(n121), .Z(n112) );
  GTECH_NOT U141 ( .A(n122), .Z(n121) );
  GTECH_AO21 U142 ( .A(n123), .B(n105), .C(n106), .Z(n120) );
  GTECH_NOT U143 ( .A(n124), .Z(n106) );
  GTECH_AO21 U144 ( .A(b[9]), .B(a[9]), .C(n125), .Z(n123) );
  GTECH_AND3 U145 ( .A(a[8]), .B(n68), .C(b[8]), .Z(n125) );
  GTECH_NAND4 U146 ( .A(n103), .B(n105), .C(n70), .D(n68), .Z(n111) );
  GTECH_XOR2 U147 ( .A(a[9]), .B(b[9]), .Z(n68) );
  GTECH_XOR2 U148 ( .A(a[8]), .B(b[8]), .Z(n70) );
  GTECH_OA21 U149 ( .A(a[10]), .B(b[10]), .C(n124), .Z(n105) );
  GTECH_NAND2 U150 ( .A(a[10]), .B(b[10]), .Z(n124) );
  GTECH_OA21 U151 ( .A(a[11]), .B(b[11]), .C(n122), .Z(n103) );
  GTECH_NAND2 U152 ( .A(a[11]), .B(b[11]), .Z(n122) );
  GTECH_AOI222 U153 ( .A(n115), .B(n126), .C(b[7]), .D(a[7]), .E(n72), .F(n127), .Z(n114) );
  GTECH_AO21 U154 ( .A(n128), .B(n75), .C(n76), .Z(n127) );
  GTECH_NOT U155 ( .A(n129), .Z(n76) );
  GTECH_AO21 U156 ( .A(b[5]), .B(a[5]), .C(n130), .Z(n128) );
  GTECH_AND3 U157 ( .A(a[4]), .B(n78), .C(b[4]), .Z(n130) );
  GTECH_AO22 U158 ( .A(b[3]), .B(a[3]), .C(n131), .D(n82), .Z(n126) );
  GTECH_XOR2 U159 ( .A(a[3]), .B(b[3]), .Z(n82) );
  GTECH_AO21 U160 ( .A(n132), .B(n85), .C(n86), .Z(n131) );
  GTECH_AND2 U161 ( .A(a[2]), .B(b[2]), .Z(n86) );
  GTECH_XOR2 U162 ( .A(a[2]), .B(b[2]), .Z(n85) );
  GTECH_AO21 U163 ( .A(b[1]), .B(a[1]), .C(n133), .Z(n132) );
  GTECH_AND3 U164 ( .A(a[0]), .B(n88), .C(b[0]), .Z(n133) );
  GTECH_XOR2 U165 ( .A(a[1]), .B(b[1]), .Z(n88) );
  GTECH_AND4 U166 ( .A(n75), .B(n80), .C(n78), .D(n72), .Z(n115) );
  GTECH_XOR2 U167 ( .A(a[7]), .B(b[7]), .Z(n72) );
  GTECH_XOR2 U168 ( .A(a[5]), .B(b[5]), .Z(n78) );
  GTECH_XOR2 U169 ( .A(a[4]), .B(b[4]), .Z(n80) );
  GTECH_OA21 U170 ( .A(a[6]), .B(b[6]), .C(n129), .Z(n75) );
  GTECH_NAND2 U171 ( .A(a[6]), .B(b[6]), .Z(n129) );
endmodule

