
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n106, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n106), .K(n106), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n243) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n106), .K(n106), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n106), .K(n106), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n106), .K(n106), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n106), .K(n106), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n106), .K(n106), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]), .QN(n260) );
  GTECH_FJK1S A_reg_15_ ( .J(n106), .K(n106), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n259) );
  GTECH_FJK1S A_reg_14_ ( .J(n106), .K(n106), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n258) );
  GTECH_FJK1S A_reg_13_ ( .J(n106), .K(n106), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n257) );
  GTECH_FJK1S A_reg_12_ ( .J(n106), .K(n106), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n256) );
  GTECH_FJK1S A_reg_11_ ( .J(n106), .K(n106), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n255) );
  GTECH_FJK1S A_reg_10_ ( .J(n106), .K(n106), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n254) );
  GTECH_FJK1S A_reg_9_ ( .J(n106), .K(n106), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n253) );
  GTECH_FJK1S A_reg_8_ ( .J(n106), .K(n106), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n252) );
  GTECH_FJK1S A_reg_7_ ( .J(n106), .K(n106), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n251) );
  GTECH_FJK1S A_reg_6_ ( .J(n106), .K(n106), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n250) );
  GTECH_FJK1S A_reg_5_ ( .J(n106), .K(n106), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n249) );
  GTECH_FJK1S A_reg_4_ ( .J(n106), .K(n106), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n248) );
  GTECH_FJK1S A_reg_3_ ( .J(n106), .K(n106), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n247) );
  GTECH_FJK1S A_reg_2_ ( .J(n106), .K(n106), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n246) );
  GTECH_FJK1S A_reg_1_ ( .J(n106), .K(n106), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n245) );
  GTECH_FJK1S A_reg_0_ ( .J(n106), .K(n106), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n244) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n106), .K(n106), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n106), .K(n106), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n106), .K(n106), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n106), .K(n106), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n106), .K(n106), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n106), .K(n106), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n106), .K(n106), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n106), .K(n106), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n106), .K(n106), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n106), .K(n106), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n106), .K(n106), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n106), .K(n106), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n106), .K(n106), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n106), .K(n106), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n106), .K(n106), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n106), .K(n106), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n106), .K(n106), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n106), .K(n106), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n106), .K(n106), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n106), .K(n106), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n106), .K(n106), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n106), .K(n106), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n106), .K(n106), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n106), .K(n106), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n106), .K(n106), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n106), .K(n106), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n106), .K(n106), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n106), .K(n106), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n106), .K(n106), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n106), .K(n106), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n106), .K(n106), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n106), .K(n106), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n106), .K(n106), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n106), .K(n106), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n106), .K(n106), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n106), .K(n106), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n106), .K(n106), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n106), .K(n106), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n106), .K(n106), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n106), .K(n106), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n106), .K(n106), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n106), .K(n106), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n106), .K(n106), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n106), .K(n106), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n106), .K(n106), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n106), .K(n106), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n106), .K(n106), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n106), .K(n106), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n106), .K(n106), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n106), .K(n106), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n106), .K(n106), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n106), .K(n106), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n106), .K(n106), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n106), .K(n106), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n106), .K(n106), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n106), .K(n106), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n106), .K(n106), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n106), .K(n106), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n106), .K(n106), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n106), .K(n106), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n106), .K(n106), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n106), .K(n106), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n106), .K(n106), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n106), .K(n106), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n106), .K(n106), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n106), .K(n106), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U245 ( .Z(n106) );
  GTECH_AND2 U246 ( .A(n261), .B(n262), .Z(N99) );
  GTECH_OAI2N2 U247 ( .A(n263), .B(n264), .C(R[15]), .D(n265), .Z(N98) );
  GTECH_OAI2N2 U248 ( .A(n13), .B(n264), .C(R[14]), .D(n265), .Z(N97) );
  GTECH_OAI2N2 U249 ( .A(n14), .B(n264), .C(R[13]), .D(n265), .Z(N96) );
  GTECH_OAI2N2 U250 ( .A(n15), .B(n264), .C(R[12]), .D(n265), .Z(N95) );
  GTECH_OAI2N2 U251 ( .A(n16), .B(n264), .C(R[11]), .D(n265), .Z(N94) );
  GTECH_OAI2N2 U252 ( .A(n17), .B(n264), .C(R[10]), .D(n265), .Z(N93) );
  GTECH_OAI2N2 U253 ( .A(n18), .B(n264), .C(R[9]), .D(n265), .Z(N92) );
  GTECH_OAI2N2 U254 ( .A(n19), .B(n264), .C(R[8]), .D(n265), .Z(N91) );
  GTECH_OAI2N2 U255 ( .A(n20), .B(n264), .C(R[7]), .D(n265), .Z(N90) );
  GTECH_OAI2N2 U256 ( .A(n21), .B(n264), .C(R[6]), .D(n265), .Z(N89) );
  GTECH_OAI2N2 U257 ( .A(n22), .B(n264), .C(R[5]), .D(n265), .Z(N88) );
  GTECH_OAI2N2 U258 ( .A(n23), .B(n264), .C(R[4]), .D(n265), .Z(N87) );
  GTECH_OAI2N2 U259 ( .A(n24), .B(n264), .C(R[3]), .D(n265), .Z(N86) );
  GTECH_OAI2N2 U260 ( .A(n25), .B(n264), .C(R[2]), .D(n265), .Z(N85) );
  GTECH_OAI2N2 U261 ( .A(n26), .B(n264), .C(R[1]), .D(n265), .Z(N84) );
  GTECH_OAI2N2 U262 ( .A(n27), .B(n264), .C(R[0]), .D(n265), .Z(N83) );
  GTECH_AND2 U263 ( .A(n261), .B(n266), .Z(N82) );
  GTECH_NOT U264 ( .A(n28), .Z(n266) );
  GTECH_AND2 U265 ( .A(M[15]), .B(n265), .Z(N42) );
  GTECH_AND2 U266 ( .A(M[14]), .B(n265), .Z(N39) );
  GTECH_AND2 U267 ( .A(M[13]), .B(n265), .Z(N38) );
  GTECH_AND2 U268 ( .A(M[12]), .B(n265), .Z(N37) );
  GTECH_AND2 U269 ( .A(M[11]), .B(n265), .Z(N36) );
  GTECH_AND2 U270 ( .A(M[10]), .B(n265), .Z(N35) );
  GTECH_AND2 U271 ( .A(M[9]), .B(n265), .Z(N34) );
  GTECH_AND2 U272 ( .A(M[8]), .B(n265), .Z(N33) );
  GTECH_AND2 U273 ( .A(M[7]), .B(n265), .Z(N32) );
  GTECH_AND2 U274 ( .A(M[6]), .B(n265), .Z(N31) );
  GTECH_AND2 U275 ( .A(M[5]), .B(n265), .Z(N30) );
  GTECH_AND2 U276 ( .A(M[4]), .B(n265), .Z(N29) );
  GTECH_AND2 U277 ( .A(M[3]), .B(n265), .Z(N28) );
  GTECH_AND2 U278 ( .A(M[2]), .B(n265), .Z(N27) );
  GTECH_AND2 U279 ( .A(M[1]), .B(n265), .Z(N26) );
  GTECH_AND2 U280 ( .A(M[0]), .B(n265), .Z(N25) );
  GTECH_OAI21 U281 ( .A(n264), .B(n267), .C(n268), .Z(N19) );
  GTECH_OR_NOT U282 ( .A(n9), .B(n269), .Z(n267) );
  GTECH_NAND3 U283 ( .A(n270), .B(n271), .C(n264), .Z(N18) );
  GTECH_AOI21 U284 ( .A(n269), .B(n272), .C(n264), .Z(N17) );
  GTECH_OR_NOT U285 ( .A(n8), .B(n273), .Z(n272) );
  GTECH_AOI21 U286 ( .A(n273), .B(n274), .C(n264), .Z(N16) );
  GTECH_OR_NOT U287 ( .A(n7), .B(n275), .Z(n274) );
  GTECH_AND2 U288 ( .A(N155), .B(n276), .Z(N152) );
  GTECH_OR_NOT U289 ( .A(N155), .B(n271), .Z(N151) );
  GTECH_AND2 U290 ( .A(N155), .B(n277), .Z(N150) );
  GTECH_MUX2 U291 ( .A(n278), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND2 U292 ( .A(n261), .B(n279), .Z(n278) );
  GTECH_AND2 U293 ( .A(N155), .B(n280), .Z(N149) );
  GTECH_AND2 U294 ( .A(N155), .B(n281), .Z(N148) );
  GTECH_AND2 U295 ( .A(N155), .B(n282), .Z(N147) );
  GTECH_AND2 U296 ( .A(N155), .B(n283), .Z(N146) );
  GTECH_AND2 U297 ( .A(N155), .B(n284), .Z(N145) );
  GTECH_AND2 U298 ( .A(N155), .B(n285), .Z(N144) );
  GTECH_AND2 U299 ( .A(N155), .B(n286), .Z(N143) );
  GTECH_AND2 U300 ( .A(N155), .B(n287), .Z(N142) );
  GTECH_AND2 U301 ( .A(N155), .B(n288), .Z(N141) );
  GTECH_AND2 U302 ( .A(N155), .B(n289), .Z(N140) );
  GTECH_NOT U303 ( .A(n290), .Z(N14) );
  GTECH_OR_NOT U304 ( .A(n279), .B(n261), .Z(n290) );
  GTECH_AND2 U305 ( .A(N155), .B(n291), .Z(N139) );
  GTECH_AND2 U306 ( .A(N155), .B(n292), .Z(N138) );
  GTECH_AND2 U307 ( .A(N155), .B(n293), .Z(N137) );
  GTECH_AND2 U308 ( .A(N155), .B(n262), .Z(N136) );
  GTECH_OAI21 U309 ( .A(n11), .B(n294), .C(n295), .Z(n262) );
  GTECH_MUX2 U310 ( .A(n296), .B(n297), .S(n298), .Z(n295) );
  GTECH_XOR2 U311 ( .A(n245), .B(n11), .Z(n298) );
  GTECH_OA22 U312 ( .A(n299), .B(n300), .C(n301), .D(n302), .Z(n297) );
  GTECH_NOT U313 ( .A(n303), .Z(n301) );
  GTECH_NOT U314 ( .A(n304), .Z(n299) );
  GTECH_OA22 U315 ( .A(n304), .B(n300), .C(n302), .D(n303), .Z(n296) );
  GTECH_AND2 U316 ( .A(N155), .B(n305), .Z(N135) );
  GTECH_NOT U317 ( .A(n263), .Z(n305) );
  GTECH_MUX2 U318 ( .A(n12), .B(n306), .S(n294), .Z(n263) );
  GTECH_AND2 U319 ( .A(n304), .B(n307), .Z(n306) );
  GTECH_OR_NOT U320 ( .A(n12), .B(n244), .Z(n307) );
  GTECH_AND2 U321 ( .A(N155), .B(n308), .Z(N134) );
  GTECH_NOT U322 ( .A(n13), .Z(n308) );
  GTECH_AND2 U323 ( .A(N155), .B(n309), .Z(N133) );
  GTECH_NOT U324 ( .A(n14), .Z(n309) );
  GTECH_AND2 U325 ( .A(N155), .B(n310), .Z(N132) );
  GTECH_NOT U326 ( .A(n15), .Z(n310) );
  GTECH_AND2 U327 ( .A(N155), .B(n311), .Z(N131) );
  GTECH_NOT U328 ( .A(n16), .Z(n311) );
  GTECH_AND2 U329 ( .A(N155), .B(n312), .Z(N130) );
  GTECH_NOT U330 ( .A(n17), .Z(n312) );
  GTECH_AND2 U331 ( .A(N155), .B(n313), .Z(N129) );
  GTECH_NOT U332 ( .A(n18), .Z(n313) );
  GTECH_AND2 U333 ( .A(N155), .B(n314), .Z(N128) );
  GTECH_NOT U334 ( .A(n19), .Z(n314) );
  GTECH_AND2 U335 ( .A(N155), .B(n315), .Z(N127) );
  GTECH_NOT U336 ( .A(n20), .Z(n315) );
  GTECH_AND2 U337 ( .A(N155), .B(n316), .Z(N126) );
  GTECH_NOT U338 ( .A(n21), .Z(n316) );
  GTECH_AND2 U339 ( .A(N155), .B(n317), .Z(N125) );
  GTECH_NOT U340 ( .A(n22), .Z(n317) );
  GTECH_AND2 U341 ( .A(N155), .B(n318), .Z(N124) );
  GTECH_NOT U342 ( .A(n23), .Z(n318) );
  GTECH_AND2 U343 ( .A(N155), .B(n319), .Z(N123) );
  GTECH_NOT U344 ( .A(n24), .Z(n319) );
  GTECH_AND2 U345 ( .A(N155), .B(n320), .Z(N122) );
  GTECH_NOT U346 ( .A(n25), .Z(n320) );
  GTECH_AND2 U347 ( .A(N155), .B(n321), .Z(N121) );
  GTECH_NOT U348 ( .A(n26), .Z(n321) );
  GTECH_AND2 U349 ( .A(N155), .B(n322), .Z(N120) );
  GTECH_NOT U350 ( .A(n27), .Z(n322) );
  GTECH_AND3 U351 ( .A(n8), .B(n7), .C(n323), .Z(N155) );
  GTECH_AND4 U352 ( .A(n279), .B(n6), .C(n271), .D(n9), .Z(n323) );
  GTECH_AND2 U353 ( .A(n261), .B(n276), .Z(N116) );
  GTECH_MUX2 U354 ( .A(n324), .B(n325), .S(n30), .Z(n276) );
  GTECH_MUX2 U355 ( .A(n326), .B(n327), .S(n260), .Z(n325) );
  GTECH_OR_NOT U356 ( .A(n328), .B(n294), .Z(n324) );
  GTECH_MUX2 U357 ( .A(n327), .B(n326), .S(n260), .Z(n328) );
  GTECH_OAI22 U358 ( .A(n302), .B(n329), .C(n330), .D(n300), .Z(n326) );
  GTECH_NOT U359 ( .A(n331), .Z(n330) );
  GTECH_NOT U360 ( .A(n332), .Z(n329) );
  GTECH_OAI22 U361 ( .A(n332), .B(n302), .C(n300), .D(n331), .Z(n327) );
  GTECH_OAI2N2 U362 ( .A(n31), .B(n333), .C(n334), .D(n335), .Z(n331) );
  GTECH_OR_NOT U363 ( .A(n259), .B(n31), .Z(n335) );
  GTECH_NOT U364 ( .A(n259), .Z(n333) );
  GTECH_ADD_ABC U365 ( .A(n31), .B(n259), .C(n336), .COUT(n332) );
  GTECH_OR_NOT U366 ( .A(N41), .B(n264), .Z(N115) );
  GTECH_OR_NOT U367 ( .A(n265), .B(n271), .Z(N41) );
  GTECH_NOT U368 ( .A(n268), .Z(n265) );
  GTECH_OR_NOT U369 ( .A(Rst), .B(Ld), .Z(n268) );
  GTECH_AND2 U370 ( .A(n261), .B(n277), .Z(N113) );
  GTECH_OAI21 U371 ( .A(n31), .B(n294), .C(n337), .Z(n277) );
  GTECH_MUX2 U372 ( .A(n338), .B(n339), .S(n340), .Z(n337) );
  GTECH_XOR2 U373 ( .A(n31), .B(n259), .Z(n340) );
  GTECH_OA22 U374 ( .A(n341), .B(n300), .C(n302), .D(n342), .Z(n339) );
  GTECH_NOT U375 ( .A(n336), .Z(n342) );
  GTECH_NOT U376 ( .A(n334), .Z(n341) );
  GTECH_OA22 U377 ( .A(n300), .B(n334), .C(n336), .D(n302), .Z(n338) );
  GTECH_ADD_ABC U378 ( .A(n32), .B(n258), .C(n343), .COUT(n336) );
  GTECH_OAI2N2 U379 ( .A(n32), .B(n344), .C(n345), .D(n346), .Z(n334) );
  GTECH_OR_NOT U380 ( .A(n258), .B(n32), .Z(n346) );
  GTECH_NOT U381 ( .A(n258), .Z(n344) );
  GTECH_AND2 U382 ( .A(n261), .B(n280), .Z(N112) );
  GTECH_OAI21 U383 ( .A(n32), .B(n294), .C(n347), .Z(n280) );
  GTECH_MUX2 U384 ( .A(n348), .B(n349), .S(n350), .Z(n347) );
  GTECH_XOR2 U385 ( .A(n32), .B(n258), .Z(n350) );
  GTECH_OA22 U386 ( .A(n351), .B(n300), .C(n302), .D(n352), .Z(n349) );
  GTECH_NOT U387 ( .A(n343), .Z(n352) );
  GTECH_NOT U388 ( .A(n345), .Z(n351) );
  GTECH_OA22 U389 ( .A(n300), .B(n345), .C(n343), .D(n302), .Z(n348) );
  GTECH_ADD_ABC U390 ( .A(n33), .B(n257), .C(n353), .COUT(n343) );
  GTECH_OAI2N2 U391 ( .A(n33), .B(n354), .C(n355), .D(n356), .Z(n345) );
  GTECH_OR_NOT U392 ( .A(n257), .B(n33), .Z(n356) );
  GTECH_NOT U393 ( .A(n257), .Z(n354) );
  GTECH_AND2 U394 ( .A(n261), .B(n281), .Z(N111) );
  GTECH_OAI21 U395 ( .A(n33), .B(n294), .C(n357), .Z(n281) );
  GTECH_MUX2 U396 ( .A(n358), .B(n359), .S(n360), .Z(n357) );
  GTECH_XOR2 U397 ( .A(n33), .B(n257), .Z(n360) );
  GTECH_OA22 U398 ( .A(n361), .B(n300), .C(n302), .D(n362), .Z(n359) );
  GTECH_NOT U399 ( .A(n353), .Z(n362) );
  GTECH_NOT U400 ( .A(n355), .Z(n361) );
  GTECH_OA22 U401 ( .A(n300), .B(n355), .C(n353), .D(n302), .Z(n358) );
  GTECH_ADD_ABC U402 ( .A(n34), .B(n256), .C(n363), .COUT(n353) );
  GTECH_OAI2N2 U403 ( .A(n34), .B(n364), .C(n365), .D(n366), .Z(n355) );
  GTECH_OR_NOT U404 ( .A(n256), .B(n34), .Z(n366) );
  GTECH_NOT U405 ( .A(n256), .Z(n364) );
  GTECH_AND2 U406 ( .A(n261), .B(n282), .Z(N110) );
  GTECH_OAI21 U407 ( .A(n34), .B(n294), .C(n367), .Z(n282) );
  GTECH_MUX2 U408 ( .A(n368), .B(n369), .S(n370), .Z(n367) );
  GTECH_XOR2 U409 ( .A(n34), .B(n256), .Z(n370) );
  GTECH_OA22 U410 ( .A(n371), .B(n300), .C(n302), .D(n372), .Z(n369) );
  GTECH_NOT U411 ( .A(n363), .Z(n372) );
  GTECH_NOT U412 ( .A(n365), .Z(n371) );
  GTECH_OA22 U413 ( .A(n300), .B(n365), .C(n363), .D(n302), .Z(n368) );
  GTECH_ADD_ABC U414 ( .A(n35), .B(n255), .C(n373), .COUT(n363) );
  GTECH_OAI2N2 U415 ( .A(n35), .B(n374), .C(n375), .D(n376), .Z(n365) );
  GTECH_OR_NOT U416 ( .A(n255), .B(n35), .Z(n376) );
  GTECH_NOT U417 ( .A(n255), .Z(n374) );
  GTECH_AND2 U418 ( .A(n261), .B(n283), .Z(N109) );
  GTECH_OAI21 U419 ( .A(n35), .B(n294), .C(n377), .Z(n283) );
  GTECH_MUX2 U420 ( .A(n378), .B(n379), .S(n380), .Z(n377) );
  GTECH_XOR2 U421 ( .A(n35), .B(n255), .Z(n380) );
  GTECH_OA22 U422 ( .A(n381), .B(n300), .C(n302), .D(n382), .Z(n379) );
  GTECH_NOT U423 ( .A(n373), .Z(n382) );
  GTECH_NOT U424 ( .A(n375), .Z(n381) );
  GTECH_OA22 U425 ( .A(n300), .B(n375), .C(n373), .D(n302), .Z(n378) );
  GTECH_ADD_ABC U426 ( .A(n36), .B(n254), .C(n383), .COUT(n373) );
  GTECH_OAI2N2 U427 ( .A(n36), .B(n384), .C(n385), .D(n386), .Z(n375) );
  GTECH_OR_NOT U428 ( .A(n254), .B(n36), .Z(n386) );
  GTECH_NOT U429 ( .A(n254), .Z(n384) );
  GTECH_AND2 U430 ( .A(n261), .B(n284), .Z(N108) );
  GTECH_OAI21 U431 ( .A(n36), .B(n294), .C(n387), .Z(n284) );
  GTECH_MUX2 U432 ( .A(n388), .B(n389), .S(n390), .Z(n387) );
  GTECH_XOR2 U433 ( .A(n36), .B(n254), .Z(n390) );
  GTECH_OA22 U434 ( .A(n391), .B(n300), .C(n302), .D(n392), .Z(n389) );
  GTECH_NOT U435 ( .A(n383), .Z(n392) );
  GTECH_NOT U436 ( .A(n385), .Z(n391) );
  GTECH_OA22 U437 ( .A(n300), .B(n385), .C(n383), .D(n302), .Z(n388) );
  GTECH_ADD_ABC U438 ( .A(n37), .B(n253), .C(n393), .COUT(n383) );
  GTECH_OAI2N2 U439 ( .A(n37), .B(n394), .C(n395), .D(n396), .Z(n385) );
  GTECH_OR_NOT U440 ( .A(n253), .B(n37), .Z(n396) );
  GTECH_NOT U441 ( .A(n253), .Z(n394) );
  GTECH_AND2 U442 ( .A(n261), .B(n285), .Z(N107) );
  GTECH_OAI21 U443 ( .A(n37), .B(n294), .C(n397), .Z(n285) );
  GTECH_MUX2 U444 ( .A(n398), .B(n399), .S(n400), .Z(n397) );
  GTECH_XOR2 U445 ( .A(n37), .B(n253), .Z(n400) );
  GTECH_OA22 U446 ( .A(n401), .B(n300), .C(n302), .D(n402), .Z(n399) );
  GTECH_NOT U447 ( .A(n393), .Z(n402) );
  GTECH_NOT U448 ( .A(n395), .Z(n401) );
  GTECH_OA22 U449 ( .A(n300), .B(n395), .C(n393), .D(n302), .Z(n398) );
  GTECH_ADD_ABC U450 ( .A(n38), .B(n252), .C(n403), .COUT(n393) );
  GTECH_OAI2N2 U451 ( .A(n38), .B(n404), .C(n405), .D(n406), .Z(n395) );
  GTECH_OR_NOT U452 ( .A(n252), .B(n38), .Z(n406) );
  GTECH_NOT U453 ( .A(n252), .Z(n404) );
  GTECH_AND2 U454 ( .A(n261), .B(n286), .Z(N106) );
  GTECH_OAI21 U455 ( .A(n38), .B(n294), .C(n407), .Z(n286) );
  GTECH_MUX2 U456 ( .A(n408), .B(n409), .S(n410), .Z(n407) );
  GTECH_XOR2 U457 ( .A(n38), .B(n252), .Z(n410) );
  GTECH_OA22 U458 ( .A(n411), .B(n300), .C(n302), .D(n412), .Z(n409) );
  GTECH_NOT U459 ( .A(n403), .Z(n412) );
  GTECH_NOT U460 ( .A(n405), .Z(n411) );
  GTECH_OA22 U461 ( .A(n300), .B(n405), .C(n403), .D(n302), .Z(n408) );
  GTECH_ADD_ABC U462 ( .A(n39), .B(n251), .C(n413), .COUT(n403) );
  GTECH_OAI2N2 U463 ( .A(n39), .B(n414), .C(n415), .D(n416), .Z(n405) );
  GTECH_OR_NOT U464 ( .A(n251), .B(n39), .Z(n416) );
  GTECH_NOT U465 ( .A(n251), .Z(n414) );
  GTECH_AND2 U466 ( .A(n261), .B(n287), .Z(N105) );
  GTECH_OAI21 U467 ( .A(n39), .B(n294), .C(n417), .Z(n287) );
  GTECH_MUX2 U468 ( .A(n418), .B(n419), .S(n420), .Z(n417) );
  GTECH_XOR2 U469 ( .A(n39), .B(n251), .Z(n420) );
  GTECH_OA22 U470 ( .A(n421), .B(n300), .C(n302), .D(n422), .Z(n419) );
  GTECH_NOT U471 ( .A(n413), .Z(n422) );
  GTECH_NOT U472 ( .A(n415), .Z(n421) );
  GTECH_OA22 U473 ( .A(n300), .B(n415), .C(n413), .D(n302), .Z(n418) );
  GTECH_ADD_ABC U474 ( .A(n40), .B(n250), .C(n423), .COUT(n413) );
  GTECH_OAI2N2 U475 ( .A(n40), .B(n424), .C(n425), .D(n426), .Z(n415) );
  GTECH_OR_NOT U476 ( .A(n250), .B(n40), .Z(n426) );
  GTECH_NOT U477 ( .A(n250), .Z(n424) );
  GTECH_AND2 U478 ( .A(n261), .B(n288), .Z(N104) );
  GTECH_OAI21 U479 ( .A(n40), .B(n294), .C(n427), .Z(n288) );
  GTECH_MUX2 U480 ( .A(n428), .B(n429), .S(n430), .Z(n427) );
  GTECH_XOR2 U481 ( .A(n40), .B(n250), .Z(n430) );
  GTECH_OA22 U482 ( .A(n431), .B(n300), .C(n302), .D(n432), .Z(n429) );
  GTECH_NOT U483 ( .A(n423), .Z(n432) );
  GTECH_NOT U484 ( .A(n425), .Z(n431) );
  GTECH_OA22 U485 ( .A(n300), .B(n425), .C(n423), .D(n302), .Z(n428) );
  GTECH_ADD_ABC U486 ( .A(n41), .B(n249), .C(n433), .COUT(n423) );
  GTECH_OAI2N2 U487 ( .A(n41), .B(n434), .C(n435), .D(n436), .Z(n425) );
  GTECH_OR_NOT U488 ( .A(n249), .B(n41), .Z(n436) );
  GTECH_NOT U489 ( .A(n249), .Z(n434) );
  GTECH_AND2 U490 ( .A(n261), .B(n289), .Z(N103) );
  GTECH_OAI21 U491 ( .A(n41), .B(n294), .C(n437), .Z(n289) );
  GTECH_MUX2 U492 ( .A(n438), .B(n439), .S(n440), .Z(n437) );
  GTECH_XOR2 U493 ( .A(n41), .B(n249), .Z(n440) );
  GTECH_OA22 U494 ( .A(n441), .B(n300), .C(n302), .D(n442), .Z(n439) );
  GTECH_NOT U495 ( .A(n433), .Z(n442) );
  GTECH_NOT U496 ( .A(n435), .Z(n441) );
  GTECH_OA22 U497 ( .A(n300), .B(n435), .C(n433), .D(n302), .Z(n438) );
  GTECH_ADD_ABC U498 ( .A(n42), .B(n248), .C(n443), .COUT(n433) );
  GTECH_OAI2N2 U499 ( .A(n42), .B(n444), .C(n445), .D(n446), .Z(n435) );
  GTECH_OR_NOT U500 ( .A(n248), .B(n42), .Z(n446) );
  GTECH_NOT U501 ( .A(n248), .Z(n444) );
  GTECH_AND2 U502 ( .A(n261), .B(n291), .Z(N102) );
  GTECH_OAI21 U503 ( .A(n42), .B(n294), .C(n447), .Z(n291) );
  GTECH_MUX2 U504 ( .A(n448), .B(n449), .S(n450), .Z(n447) );
  GTECH_XOR2 U505 ( .A(n42), .B(n248), .Z(n450) );
  GTECH_OA22 U506 ( .A(n451), .B(n300), .C(n302), .D(n452), .Z(n449) );
  GTECH_NOT U507 ( .A(n443), .Z(n452) );
  GTECH_NOT U508 ( .A(n445), .Z(n451) );
  GTECH_OA22 U509 ( .A(n300), .B(n445), .C(n443), .D(n302), .Z(n448) );
  GTECH_ADD_ABC U510 ( .A(n43), .B(n247), .C(n453), .COUT(n443) );
  GTECH_OAI2N2 U511 ( .A(n43), .B(n454), .C(n455), .D(n456), .Z(n445) );
  GTECH_OR_NOT U512 ( .A(n247), .B(n43), .Z(n456) );
  GTECH_NOT U513 ( .A(n247), .Z(n454) );
  GTECH_AND2 U514 ( .A(n261), .B(n292), .Z(N101) );
  GTECH_OAI21 U515 ( .A(n43), .B(n294), .C(n457), .Z(n292) );
  GTECH_MUX2 U516 ( .A(n458), .B(n459), .S(n460), .Z(n457) );
  GTECH_XOR2 U517 ( .A(n43), .B(n247), .Z(n460) );
  GTECH_OA22 U518 ( .A(n461), .B(n300), .C(n302), .D(n462), .Z(n459) );
  GTECH_NOT U519 ( .A(n453), .Z(n462) );
  GTECH_NOT U520 ( .A(n455), .Z(n461) );
  GTECH_OA22 U521 ( .A(n300), .B(n455), .C(n453), .D(n302), .Z(n458) );
  GTECH_ADD_ABC U522 ( .A(n29), .B(n246), .C(n463), .COUT(n453) );
  GTECH_OAI2N2 U523 ( .A(n29), .B(n464), .C(n465), .D(n466), .Z(n455) );
  GTECH_OR_NOT U524 ( .A(n246), .B(n29), .Z(n466) );
  GTECH_NOT U525 ( .A(n246), .Z(n464) );
  GTECH_AND2 U526 ( .A(n261), .B(n293), .Z(N100) );
  GTECH_OAI21 U527 ( .A(n29), .B(n294), .C(n467), .Z(n293) );
  GTECH_MUX2 U528 ( .A(n468), .B(n469), .S(n470), .Z(n467) );
  GTECH_XOR2 U529 ( .A(n29), .B(n246), .Z(n470) );
  GTECH_OA22 U530 ( .A(n471), .B(n300), .C(n302), .D(n472), .Z(n469) );
  GTECH_NOT U531 ( .A(n463), .Z(n472) );
  GTECH_NOT U532 ( .A(n465), .Z(n471) );
  GTECH_OA22 U533 ( .A(n300), .B(n465), .C(n463), .D(n302), .Z(n468) );
  GTECH_ADD_ABC U534 ( .A(n245), .B(n11), .C(n303), .COUT(n463) );
  GTECH_OR_NOT U535 ( .A(n244), .B(n473), .Z(n303) );
  GTECH_NOT U536 ( .A(n12), .Z(n473) );
  GTECH_OAI2N2 U537 ( .A(n11), .B(n474), .C(n304), .D(n475), .Z(n465) );
  GTECH_OR_NOT U538 ( .A(n245), .B(n11), .Z(n475) );
  GTECH_OR_NOT U539 ( .A(n244), .B(n12), .Z(n304) );
  GTECH_NOT U540 ( .A(n245), .Z(n474) );
  GTECH_OR_NOT U541 ( .A(n476), .B(n302), .Z(n294) );
  GTECH_OR_NOT U542 ( .A(n10), .B(n28), .Z(n302) );
  GTECH_NOT U543 ( .A(n300), .Z(n476) );
  GTECH_OR_NOT U544 ( .A(n28), .B(n10), .Z(n300) );
  GTECH_NOT U545 ( .A(n264), .Z(n261) );
  GTECH_NAND3 U546 ( .A(n270), .B(n271), .C(n477), .Z(n264) );
  GTECH_OR_NOT U547 ( .A(n269), .B(n9), .Z(n477) );
  GTECH_OR_NOT U548 ( .A(n273), .B(n8), .Z(n269) );
  GTECH_OR_NOT U549 ( .A(n275), .B(n7), .Z(n273) );
  GTECH_OR_NOT U550 ( .A(n279), .B(n6), .Z(n275) );
  GTECH_NOT U551 ( .A(n243), .Z(n279) );
  GTECH_NOT U552 ( .A(Rst), .Z(n271) );
  GTECH_NOT U553 ( .A(Ld), .Z(n270) );
endmodule

