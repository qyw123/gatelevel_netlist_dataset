
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143;

  GTECH_XNOR2 U92 ( .A(n73), .B(n74), .Z(sum[9]) );
  GTECH_XOR2 U93 ( .A(n75), .B(n76), .Z(sum[8]) );
  GTECH_XOR2 U94 ( .A(n77), .B(n78), .Z(sum[7]) );
  GTECH_OAI21 U95 ( .A(n79), .B(n80), .C(n81), .Z(n78) );
  GTECH_XOR2 U96 ( .A(n79), .B(n80), .Z(sum[6]) );
  GTECH_NOT U97 ( .A(n82), .Z(n80) );
  GTECH_OAI21 U98 ( .A(n83), .B(n84), .C(n85), .Z(n82) );
  GTECH_XOR2 U99 ( .A(n83), .B(n84), .Z(sum[5]) );
  GTECH_AOI22 U100 ( .A(b[4]), .B(a[4]), .C(n86), .D(n87), .Z(n83) );
  GTECH_XOR2 U101 ( .A(n87), .B(n86), .Z(sum[4]) );
  GTECH_XNOR2 U102 ( .A(n88), .B(n89), .Z(sum[3]) );
  GTECH_AOI21 U103 ( .A(n90), .B(n91), .C(n92), .Z(n89) );
  GTECH_XOR2 U104 ( .A(n90), .B(n91), .Z(sum[2]) );
  GTECH_AO22 U105 ( .A(n93), .B(n94), .C(b[1]), .D(a[1]), .Z(n91) );
  GTECH_XOR2 U106 ( .A(n94), .B(n93), .Z(sum[1]) );
  GTECH_AO22 U107 ( .A(n95), .B(cin), .C(a[0]), .D(b[0]), .Z(n93) );
  GTECH_XOR2 U108 ( .A(n96), .B(n97), .Z(sum[15]) );
  GTECH_AOI21 U109 ( .A(n98), .B(n99), .C(n100), .Z(n97) );
  GTECH_XNOR2 U110 ( .A(n99), .B(n101), .Z(sum[14]) );
  GTECH_OAI21 U111 ( .A(n102), .B(n103), .C(n104), .Z(n99) );
  GTECH_XOR2 U112 ( .A(n103), .B(n102), .Z(sum[13]) );
  GTECH_AOI21 U113 ( .A(cout), .B(n105), .C(n106), .Z(n102) );
  GTECH_NOT U114 ( .A(n107), .Z(n106) );
  GTECH_XOR2 U115 ( .A(cout), .B(n105), .Z(sum[12]) );
  GTECH_NOT U116 ( .A(n108), .Z(n105) );
  GTECH_XOR2 U117 ( .A(n109), .B(n110), .Z(sum[11]) );
  GTECH_AOI21 U118 ( .A(n111), .B(n112), .C(n113), .Z(n110) );
  GTECH_XNOR2 U119 ( .A(n112), .B(n114), .Z(sum[10]) );
  GTECH_OAI2N2 U120 ( .A(n115), .B(n73), .C(b[9]), .D(a[9]), .Z(n112) );
  GTECH_NOT U121 ( .A(n74), .Z(n115) );
  GTECH_OAI21 U122 ( .A(n75), .B(n76), .C(n116), .Z(n74) );
  GTECH_NOT U123 ( .A(n117), .Z(n75) );
  GTECH_XOR2 U124 ( .A(cin), .B(n95), .Z(sum[0]) );
  GTECH_AO21 U125 ( .A(n117), .B(n118), .C(n119), .Z(cout) );
  GTECH_AO21 U126 ( .A(n86), .B(n120), .C(n121), .Z(n117) );
  GTECH_AO21 U127 ( .A(n122), .B(cin), .C(n123), .Z(n86) );
  GTECH_NOT U128 ( .A(n124), .Z(Pm) );
  GTECH_NAND3 U129 ( .A(n118), .B(n122), .C(n120), .Z(n124) );
  GTECH_AND5 U130 ( .A(n90), .B(n94), .C(n88), .D(n125), .E(n95), .Z(n122) );
  GTECH_XOR2 U131 ( .A(a[0]), .B(b[0]), .Z(n95) );
  GTECH_AO21 U132 ( .A(n126), .B(n118), .C(n119), .Z(Gm) );
  GTECH_OAI2N2 U133 ( .A(n127), .B(n96), .C(b[15]), .D(a[15]), .Z(n119) );
  GTECH_AOI21 U134 ( .A(n98), .B(n128), .C(n100), .Z(n127) );
  GTECH_NOT U135 ( .A(n129), .Z(n100) );
  GTECH_OAI21 U136 ( .A(n107), .B(n103), .C(n104), .Z(n128) );
  GTECH_NOT U137 ( .A(n101), .Z(n98) );
  GTECH_NOR4 U138 ( .A(n108), .B(n101), .C(n103), .D(n96), .Z(n118) );
  GTECH_XNOR2 U139 ( .A(a[15]), .B(b[15]), .Z(n96) );
  GTECH_OAI21 U140 ( .A(b[13]), .B(a[13]), .C(n104), .Z(n103) );
  GTECH_NAND2 U141 ( .A(a[13]), .B(b[13]), .Z(n104) );
  GTECH_OAI21 U142 ( .A(b[14]), .B(a[14]), .C(n129), .Z(n101) );
  GTECH_NAND2 U143 ( .A(a[14]), .B(b[14]), .Z(n129) );
  GTECH_OAI21 U144 ( .A(b[12]), .B(a[12]), .C(n107), .Z(n108) );
  GTECH_NAND2 U145 ( .A(b[12]), .B(a[12]), .Z(n107) );
  GTECH_AO21 U146 ( .A(n120), .B(n123), .C(n121), .Z(n126) );
  GTECH_OAI2N2 U147 ( .A(n130), .B(n109), .C(b[11]), .D(a[11]), .Z(n121) );
  GTECH_AOI21 U148 ( .A(n111), .B(n131), .C(n113), .Z(n130) );
  GTECH_NOT U149 ( .A(n132), .Z(n113) );
  GTECH_OAI2N2 U150 ( .A(n73), .B(n116), .C(b[9]), .D(a[9]), .Z(n131) );
  GTECH_NOT U151 ( .A(n114), .Z(n111) );
  GTECH_NOT U152 ( .A(n133), .Z(n123) );
  GTECH_AOI222 U153 ( .A(a[7]), .B(b[7]), .C(n125), .D(n134), .E(n77), .F(n135), .Z(n133) );
  GTECH_NAND2 U154 ( .A(n136), .B(n81), .Z(n135) );
  GTECH_NAND2 U155 ( .A(a[6]), .B(b[6]), .Z(n81) );
  GTECH_AO21 U156 ( .A(n137), .B(n85), .C(n79), .Z(n136) );
  GTECH_NOT U157 ( .A(n138), .Z(n79) );
  GTECH_NAND3 U158 ( .A(n139), .B(b[4]), .C(a[4]), .Z(n137) );
  GTECH_AO22 U159 ( .A(n140), .B(n88), .C(b[3]), .D(a[3]), .Z(n134) );
  GTECH_XOR2 U160 ( .A(a[3]), .B(b[3]), .Z(n88) );
  GTECH_AO21 U161 ( .A(n90), .B(n141), .C(n92), .Z(n140) );
  GTECH_AND2 U162 ( .A(a[2]), .B(b[2]), .Z(n92) );
  GTECH_AO21 U163 ( .A(b[1]), .B(a[1]), .C(n142), .Z(n141) );
  GTECH_NOT U164 ( .A(n143), .Z(n142) );
  GTECH_NAND3 U165 ( .A(a[0]), .B(n94), .C(b[0]), .Z(n143) );
  GTECH_XOR2 U166 ( .A(a[1]), .B(b[1]), .Z(n94) );
  GTECH_XOR2 U167 ( .A(a[2]), .B(b[2]), .Z(n90) );
  GTECH_AND4 U168 ( .A(n139), .B(n87), .C(n138), .D(n77), .Z(n125) );
  GTECH_XOR2 U169 ( .A(a[7]), .B(b[7]), .Z(n77) );
  GTECH_XOR2 U170 ( .A(a[6]), .B(b[6]), .Z(n138) );
  GTECH_XOR2 U171 ( .A(a[4]), .B(b[4]), .Z(n87) );
  GTECH_NOT U172 ( .A(n84), .Z(n139) );
  GTECH_OAI21 U173 ( .A(b[5]), .B(a[5]), .C(n85), .Z(n84) );
  GTECH_NAND2 U174 ( .A(b[5]), .B(a[5]), .Z(n85) );
  GTECH_NOR4 U175 ( .A(n76), .B(n114), .C(n109), .D(n73), .Z(n120) );
  GTECH_XNOR2 U176 ( .A(a[9]), .B(b[9]), .Z(n73) );
  GTECH_XNOR2 U177 ( .A(a[11]), .B(b[11]), .Z(n109) );
  GTECH_OAI21 U178 ( .A(b[10]), .B(a[10]), .C(n132), .Z(n114) );
  GTECH_NAND2 U179 ( .A(a[10]), .B(b[10]), .Z(n132) );
  GTECH_OAI21 U180 ( .A(b[8]), .B(a[8]), .C(n116), .Z(n76) );
  GTECH_NAND2 U181 ( .A(b[8]), .B(a[8]), .Z(n116) );
endmodule

