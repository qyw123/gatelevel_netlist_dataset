
module counter10 ( clk, reset, q );
  output [3:0] q;
  input clk, reset;
  wire   N7, N8, N9, N10, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29;

  GTECH_FD1 q_reg_0_ ( .D(N7), .CP(clk), .Q(q[0]) );
  GTECH_FD1 q_reg_3_ ( .D(N10), .CP(clk), .Q(q[3]) );
  GTECH_FD1 q_reg_1_ ( .D(N8), .CP(clk), .Q(q[1]) );
  GTECH_FD1 q_reg_2_ ( .D(N9), .CP(clk), .Q(q[2]) );
  GTECH_NOR3 U16 ( .A(n19), .B(reset), .C(q[3]), .Z(N9) );
  GTECH_XOR2 U17 ( .A(n20), .B(q[2]), .Z(n19) );
  GTECH_AND4 U18 ( .A(n21), .B(n20), .C(n22), .D(n23), .Z(N8) );
  GTECH_NOT U19 ( .A(reset), .Z(n23) );
  GTECH_NOT U20 ( .A(q[3]), .Z(n22) );
  GTECH_NOR3 U21 ( .A(n24), .B(reset), .C(q[0]), .Z(N7) );
  GTECH_OA21 U22 ( .A(q[2]), .B(q[1]), .C(q[3]), .Z(n24) );
  GTECH_NOR3 U23 ( .A(n25), .B(n26), .C(n27), .Z(N10) );
  GTECH_OA21 U24 ( .A(n20), .B(q[3]), .C(q[2]), .Z(n27) );
  GTECH_AO21 U25 ( .A(n21), .B(n20), .C(reset), .Z(n26) );
  GTECH_NAND2 U26 ( .A(n28), .B(n29), .Z(n21) );
  GTECH_NOT U27 ( .A(q[0]), .Z(n29) );
  GTECH_NOT U28 ( .A(q[1]), .Z(n28) );
  GTECH_AOI21 U29 ( .A(n20), .B(q[3]), .C(q[2]), .Z(n25) );
  GTECH_NAND2 U30 ( .A(q[1]), .B(q[0]), .Z(n20) );
endmodule

