
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n105, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n105), .K(n105), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n242) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n105), .K(n105), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n105), .K(n105), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n105), .K(n105), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n105), .K(n105), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n105), .K(n105), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]), .QN(n259) );
  GTECH_FJK1S A_reg_15_ ( .J(n105), .K(n105), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n258) );
  GTECH_FJK1S A_reg_14_ ( .J(n105), .K(n105), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n257) );
  GTECH_FJK1S A_reg_13_ ( .J(n105), .K(n105), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n256) );
  GTECH_FJK1S A_reg_12_ ( .J(n105), .K(n105), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n255) );
  GTECH_FJK1S A_reg_11_ ( .J(n105), .K(n105), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n254) );
  GTECH_FJK1S A_reg_10_ ( .J(n105), .K(n105), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n253) );
  GTECH_FJK1S A_reg_9_ ( .J(n105), .K(n105), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n252) );
  GTECH_FJK1S A_reg_8_ ( .J(n105), .K(n105), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n251) );
  GTECH_FJK1S A_reg_7_ ( .J(n105), .K(n105), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n250) );
  GTECH_FJK1S A_reg_6_ ( .J(n105), .K(n105), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n249) );
  GTECH_FJK1S A_reg_5_ ( .J(n105), .K(n105), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n248) );
  GTECH_FJK1S A_reg_4_ ( .J(n105), .K(n105), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n247) );
  GTECH_FJK1S A_reg_3_ ( .J(n105), .K(n105), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n246) );
  GTECH_FJK1S A_reg_2_ ( .J(n105), .K(n105), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n245) );
  GTECH_FJK1S A_reg_1_ ( .J(n105), .K(n105), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n244) );
  GTECH_FJK1S A_reg_0_ ( .J(n105), .K(n105), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n243) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n105), .K(n105), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n105), .K(n105), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n105), .K(n105), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n105), .K(n105), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n105), .K(n105), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n105), .K(n105), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n105), .K(n105), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n105), .K(n105), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n105), .K(n105), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n105), .K(n105), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n105), .K(n105), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n105), .K(n105), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n105), .K(n105), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n105), .K(n105), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n105), .K(n105), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n105), .K(n105), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n105), .K(n105), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n105), .K(n105), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n105), .K(n105), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n105), .K(n105), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n105), .K(n105), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n105), .K(n105), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n105), .K(n105), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n105), .K(n105), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n105), .K(n105), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n105), .K(n105), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n105), .K(n105), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n105), .K(n105), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n105), .K(n105), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n105), .K(n105), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n105), .K(n105), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n105), .K(n105), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n105), .K(n105), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n105), .K(n105), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n105), .K(n105), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n105), .K(n105), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n105), .K(n105), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n105), .K(n105), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n105), .K(n105), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n105), .K(n105), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n105), .K(n105), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n105), .K(n105), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n105), .K(n105), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n105), .K(n105), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n105), .K(n105), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n105), .K(n105), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n105), .K(n105), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n105), .K(n105), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n105), .K(n105), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n105), .K(n105), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n105), .K(n105), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n105), .K(n105), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n105), .K(n105), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n105), .K(n105), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n105), .K(n105), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n105), .K(n105), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n105), .K(n105), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n105), .K(n105), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n105), .K(n105), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n105), .K(n105), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n105), .K(n105), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n105), .K(n105), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n105), .K(n105), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n105), .K(n105), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n105), .K(n105), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n105), .K(n105), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U244 ( .Z(n105) );
  GTECH_AND2 U245 ( .A(n260), .B(n261), .Z(N99) );
  GTECH_OAI2N2 U246 ( .A(n262), .B(n263), .C(R[15]), .D(n264), .Z(N98) );
  GTECH_OAI2N2 U247 ( .A(n13), .B(n263), .C(R[14]), .D(n264), .Z(N97) );
  GTECH_OAI2N2 U248 ( .A(n14), .B(n263), .C(R[13]), .D(n264), .Z(N96) );
  GTECH_OAI2N2 U249 ( .A(n15), .B(n263), .C(R[12]), .D(n264), .Z(N95) );
  GTECH_OAI2N2 U250 ( .A(n16), .B(n263), .C(R[11]), .D(n264), .Z(N94) );
  GTECH_OAI2N2 U251 ( .A(n17), .B(n263), .C(R[10]), .D(n264), .Z(N93) );
  GTECH_OAI2N2 U252 ( .A(n18), .B(n263), .C(R[9]), .D(n264), .Z(N92) );
  GTECH_OAI2N2 U253 ( .A(n19), .B(n263), .C(R[8]), .D(n264), .Z(N91) );
  GTECH_OAI2N2 U254 ( .A(n20), .B(n263), .C(R[7]), .D(n264), .Z(N90) );
  GTECH_OAI2N2 U255 ( .A(n21), .B(n263), .C(R[6]), .D(n264), .Z(N89) );
  GTECH_OAI2N2 U256 ( .A(n22), .B(n263), .C(R[5]), .D(n264), .Z(N88) );
  GTECH_OAI2N2 U257 ( .A(n23), .B(n263), .C(R[4]), .D(n264), .Z(N87) );
  GTECH_OAI2N2 U258 ( .A(n24), .B(n263), .C(R[3]), .D(n264), .Z(N86) );
  GTECH_OAI2N2 U259 ( .A(n25), .B(n263), .C(R[2]), .D(n264), .Z(N85) );
  GTECH_OAI2N2 U260 ( .A(n26), .B(n263), .C(R[1]), .D(n264), .Z(N84) );
  GTECH_OAI2N2 U261 ( .A(n27), .B(n263), .C(R[0]), .D(n264), .Z(N83) );
  GTECH_AND2 U262 ( .A(n260), .B(n265), .Z(N82) );
  GTECH_AND2 U263 ( .A(M[15]), .B(n264), .Z(N42) );
  GTECH_AND2 U264 ( .A(M[14]), .B(n264), .Z(N39) );
  GTECH_AND2 U265 ( .A(M[13]), .B(n264), .Z(N38) );
  GTECH_AND2 U266 ( .A(M[12]), .B(n264), .Z(N37) );
  GTECH_AND2 U267 ( .A(M[11]), .B(n264), .Z(N36) );
  GTECH_AND2 U268 ( .A(M[10]), .B(n264), .Z(N35) );
  GTECH_AND2 U269 ( .A(M[9]), .B(n264), .Z(N34) );
  GTECH_AND2 U270 ( .A(M[8]), .B(n264), .Z(N33) );
  GTECH_AND2 U271 ( .A(M[7]), .B(n264), .Z(N32) );
  GTECH_AND2 U272 ( .A(M[6]), .B(n264), .Z(N31) );
  GTECH_AND2 U273 ( .A(M[5]), .B(n264), .Z(N30) );
  GTECH_AND2 U274 ( .A(M[4]), .B(n264), .Z(N29) );
  GTECH_AND2 U275 ( .A(M[3]), .B(n264), .Z(N28) );
  GTECH_AND2 U276 ( .A(M[2]), .B(n264), .Z(N27) );
  GTECH_AND2 U277 ( .A(M[1]), .B(n264), .Z(N26) );
  GTECH_AND2 U278 ( .A(M[0]), .B(n264), .Z(N25) );
  GTECH_NOT U279 ( .A(n266), .Z(n264) );
  GTECH_NAND2 U280 ( .A(n266), .B(n267), .Z(N19) );
  GTECH_NAND3 U281 ( .A(n268), .B(n269), .C(n260), .Z(n267) );
  GTECH_NAND2 U282 ( .A(n270), .B(n263), .Z(N18) );
  GTECH_AND2 U283 ( .A(n260), .B(n271), .Z(N17) );
  GTECH_OAI21 U284 ( .A(n8), .B(n272), .C(n268), .Z(n271) );
  GTECH_AND2 U285 ( .A(n260), .B(n273), .Z(N16) );
  GTECH_OAI21 U286 ( .A(n7), .B(n274), .C(n275), .Z(n273) );
  GTECH_AND2 U287 ( .A(N155), .B(n276), .Z(N152) );
  GTECH_NAND2 U288 ( .A(n277), .B(n278), .Z(N151) );
  GTECH_AND2 U289 ( .A(N155), .B(n279), .Z(N150) );
  GTECH_MUX2 U290 ( .A(n280), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND2 U291 ( .A(n260), .B(n281), .Z(n280) );
  GTECH_AND2 U292 ( .A(N155), .B(n282), .Z(N149) );
  GTECH_AND2 U293 ( .A(N155), .B(n283), .Z(N148) );
  GTECH_AND2 U294 ( .A(N155), .B(n284), .Z(N147) );
  GTECH_AND2 U295 ( .A(N155), .B(n285), .Z(N146) );
  GTECH_AND2 U296 ( .A(N155), .B(n286), .Z(N145) );
  GTECH_AND2 U297 ( .A(N155), .B(n287), .Z(N144) );
  GTECH_AND2 U298 ( .A(N155), .B(n288), .Z(N143) );
  GTECH_AND2 U299 ( .A(N155), .B(n289), .Z(N142) );
  GTECH_AND2 U300 ( .A(N155), .B(n290), .Z(N141) );
  GTECH_AND2 U301 ( .A(N155), .B(n291), .Z(N140) );
  GTECH_NOT U302 ( .A(n292), .Z(N14) );
  GTECH_NAND2 U303 ( .A(n260), .B(n242), .Z(n292) );
  GTECH_AND2 U304 ( .A(N155), .B(n293), .Z(N139) );
  GTECH_AND2 U305 ( .A(N155), .B(n294), .Z(N138) );
  GTECH_AND2 U306 ( .A(N155), .B(n295), .Z(N137) );
  GTECH_AND2 U307 ( .A(N155), .B(n261), .Z(N136) );
  GTECH_OAI21 U308 ( .A(n11), .B(n296), .C(n297), .Z(n261) );
  GTECH_MUX2 U309 ( .A(n298), .B(n299), .S(n300), .Z(n297) );
  GTECH_XOR2 U310 ( .A(n244), .B(n11), .Z(n300) );
  GTECH_OA22 U311 ( .A(n301), .B(n302), .C(n303), .D(n304), .Z(n299) );
  GTECH_OA22 U312 ( .A(n302), .B(n305), .C(n304), .D(n306), .Z(n298) );
  GTECH_AND2 U313 ( .A(N155), .B(n307), .Z(N135) );
  GTECH_NOT U314 ( .A(n262), .Z(n307) );
  GTECH_MUX2 U315 ( .A(n12), .B(n308), .S(n296), .Z(n262) );
  GTECH_OA21 U316 ( .A(n309), .B(n12), .C(n305), .Z(n308) );
  GTECH_AND2 U317 ( .A(N155), .B(n310), .Z(N134) );
  GTECH_NOT U318 ( .A(n13), .Z(n310) );
  GTECH_AND2 U319 ( .A(N155), .B(n311), .Z(N133) );
  GTECH_NOT U320 ( .A(n14), .Z(n311) );
  GTECH_AND2 U321 ( .A(N155), .B(n312), .Z(N132) );
  GTECH_NOT U322 ( .A(n15), .Z(n312) );
  GTECH_AND2 U323 ( .A(N155), .B(n313), .Z(N131) );
  GTECH_NOT U324 ( .A(n16), .Z(n313) );
  GTECH_AND2 U325 ( .A(N155), .B(n314), .Z(N130) );
  GTECH_NOT U326 ( .A(n17), .Z(n314) );
  GTECH_AND2 U327 ( .A(N155), .B(n315), .Z(N129) );
  GTECH_NOT U328 ( .A(n18), .Z(n315) );
  GTECH_AND2 U329 ( .A(N155), .B(n316), .Z(N128) );
  GTECH_NOT U330 ( .A(n19), .Z(n316) );
  GTECH_AND2 U331 ( .A(N155), .B(n317), .Z(N127) );
  GTECH_NOT U332 ( .A(n20), .Z(n317) );
  GTECH_AND2 U333 ( .A(N155), .B(n318), .Z(N126) );
  GTECH_NOT U334 ( .A(n21), .Z(n318) );
  GTECH_AND2 U335 ( .A(N155), .B(n319), .Z(N125) );
  GTECH_NOT U336 ( .A(n22), .Z(n319) );
  GTECH_AND2 U337 ( .A(N155), .B(n320), .Z(N124) );
  GTECH_NOT U338 ( .A(n23), .Z(n320) );
  GTECH_AND2 U339 ( .A(N155), .B(n321), .Z(N123) );
  GTECH_NOT U340 ( .A(n24), .Z(n321) );
  GTECH_AND2 U341 ( .A(N155), .B(n322), .Z(N122) );
  GTECH_NOT U342 ( .A(n25), .Z(n322) );
  GTECH_AND2 U343 ( .A(N155), .B(n323), .Z(N121) );
  GTECH_NOT U344 ( .A(n26), .Z(n323) );
  GTECH_AND2 U345 ( .A(N155), .B(n324), .Z(N120) );
  GTECH_NOT U346 ( .A(n27), .Z(n324) );
  GTECH_NOT U347 ( .A(n278), .Z(N155) );
  GTECH_NAND4 U348 ( .A(n8), .B(n7), .C(n9), .D(n325), .Z(n278) );
  GTECH_AND3 U349 ( .A(n277), .B(n281), .C(n6), .Z(n325) );
  GTECH_NOT U350 ( .A(n242), .Z(n281) );
  GTECH_AND2 U351 ( .A(n260), .B(n276), .Z(N116) );
  GTECH_MUX2 U352 ( .A(n326), .B(n327), .S(n30), .Z(n276) );
  GTECH_MUX2 U353 ( .A(n328), .B(n329), .S(n259), .Z(n327) );
  GTECH_NAND2 U354 ( .A(n330), .B(n296), .Z(n326) );
  GTECH_MUX2 U355 ( .A(n331), .B(n332), .S(n259), .Z(n330) );
  GTECH_NOT U356 ( .A(n328), .Z(n332) );
  GTECH_OAI22 U357 ( .A(n304), .B(n333), .C(n302), .D(n334), .Z(n328) );
  GTECH_NOT U358 ( .A(n329), .Z(n331) );
  GTECH_OAI22 U359 ( .A(n335), .B(n304), .C(n336), .D(n302), .Z(n329) );
  GTECH_NOT U360 ( .A(n334), .Z(n336) );
  GTECH_OAI21 U361 ( .A(n258), .B(n337), .C(n338), .Z(n334) );
  GTECH_OAI21 U362 ( .A(n31), .B(n339), .C(n340), .Z(n338) );
  GTECH_NOT U363 ( .A(n333), .Z(n335) );
  GTECH_OAI21 U364 ( .A(n31), .B(n258), .C(n341), .Z(n333) );
  GTECH_OAI21 U365 ( .A(n339), .B(n337), .C(n342), .Z(n341) );
  GTECH_NOT U366 ( .A(n31), .Z(n337) );
  GTECH_NOT U367 ( .A(n258), .Z(n339) );
  GTECH_NAND2 U368 ( .A(n263), .B(n343), .Z(N115) );
  GTECH_NOT U369 ( .A(N41), .Z(n343) );
  GTECH_NAND2 U370 ( .A(n277), .B(n266), .Z(N41) );
  GTECH_NAND2 U371 ( .A(Ld), .B(n277), .Z(n266) );
  GTECH_AND2 U372 ( .A(n260), .B(n279), .Z(N113) );
  GTECH_MUX2 U373 ( .A(n344), .B(n345), .S(n31), .Z(n279) );
  GTECH_MUX2 U374 ( .A(n346), .B(n347), .S(n258), .Z(n345) );
  GTECH_NAND2 U375 ( .A(n348), .B(n296), .Z(n344) );
  GTECH_MUX2 U376 ( .A(n349), .B(n350), .S(n258), .Z(n348) );
  GTECH_NOT U377 ( .A(n346), .Z(n350) );
  GTECH_OAI22 U378 ( .A(n304), .B(n342), .C(n302), .D(n340), .Z(n346) );
  GTECH_NOT U379 ( .A(n347), .Z(n349) );
  GTECH_OAI22 U380 ( .A(n351), .B(n304), .C(n352), .D(n302), .Z(n347) );
  GTECH_NOT U381 ( .A(n340), .Z(n352) );
  GTECH_OAI21 U382 ( .A(n257), .B(n353), .C(n354), .Z(n340) );
  GTECH_OAI21 U383 ( .A(n32), .B(n355), .C(n356), .Z(n354) );
  GTECH_NOT U384 ( .A(n342), .Z(n351) );
  GTECH_OAI21 U385 ( .A(n32), .B(n257), .C(n357), .Z(n342) );
  GTECH_OAI21 U386 ( .A(n355), .B(n353), .C(n358), .Z(n357) );
  GTECH_NOT U387 ( .A(n32), .Z(n353) );
  GTECH_NOT U388 ( .A(n257), .Z(n355) );
  GTECH_AND2 U389 ( .A(n260), .B(n282), .Z(N112) );
  GTECH_MUX2 U390 ( .A(n359), .B(n360), .S(n32), .Z(n282) );
  GTECH_MUX2 U391 ( .A(n361), .B(n362), .S(n257), .Z(n360) );
  GTECH_NAND2 U392 ( .A(n363), .B(n296), .Z(n359) );
  GTECH_MUX2 U393 ( .A(n364), .B(n365), .S(n257), .Z(n363) );
  GTECH_NOT U394 ( .A(n361), .Z(n365) );
  GTECH_OAI22 U395 ( .A(n304), .B(n358), .C(n302), .D(n356), .Z(n361) );
  GTECH_NOT U396 ( .A(n362), .Z(n364) );
  GTECH_OAI22 U397 ( .A(n366), .B(n304), .C(n367), .D(n302), .Z(n362) );
  GTECH_NOT U398 ( .A(n356), .Z(n367) );
  GTECH_OAI21 U399 ( .A(n256), .B(n368), .C(n369), .Z(n356) );
  GTECH_OAI21 U400 ( .A(n33), .B(n370), .C(n371), .Z(n369) );
  GTECH_NOT U401 ( .A(n358), .Z(n366) );
  GTECH_OAI21 U402 ( .A(n33), .B(n256), .C(n372), .Z(n358) );
  GTECH_OAI21 U403 ( .A(n370), .B(n368), .C(n373), .Z(n372) );
  GTECH_NOT U404 ( .A(n33), .Z(n368) );
  GTECH_NOT U405 ( .A(n256), .Z(n370) );
  GTECH_AND2 U406 ( .A(n260), .B(n283), .Z(N111) );
  GTECH_MUX2 U407 ( .A(n374), .B(n375), .S(n33), .Z(n283) );
  GTECH_MUX2 U408 ( .A(n376), .B(n377), .S(n256), .Z(n375) );
  GTECH_NAND2 U409 ( .A(n378), .B(n296), .Z(n374) );
  GTECH_MUX2 U410 ( .A(n379), .B(n380), .S(n256), .Z(n378) );
  GTECH_NOT U411 ( .A(n376), .Z(n380) );
  GTECH_OAI22 U412 ( .A(n304), .B(n373), .C(n302), .D(n371), .Z(n376) );
  GTECH_NOT U413 ( .A(n377), .Z(n379) );
  GTECH_OAI22 U414 ( .A(n381), .B(n304), .C(n382), .D(n302), .Z(n377) );
  GTECH_NOT U415 ( .A(n371), .Z(n382) );
  GTECH_OAI21 U416 ( .A(n255), .B(n383), .C(n384), .Z(n371) );
  GTECH_OAI21 U417 ( .A(n34), .B(n385), .C(n386), .Z(n384) );
  GTECH_NOT U418 ( .A(n373), .Z(n381) );
  GTECH_OAI21 U419 ( .A(n34), .B(n255), .C(n387), .Z(n373) );
  GTECH_OAI21 U420 ( .A(n385), .B(n383), .C(n388), .Z(n387) );
  GTECH_NOT U421 ( .A(n34), .Z(n383) );
  GTECH_NOT U422 ( .A(n255), .Z(n385) );
  GTECH_AND2 U423 ( .A(n260), .B(n284), .Z(N110) );
  GTECH_MUX2 U424 ( .A(n389), .B(n390), .S(n34), .Z(n284) );
  GTECH_MUX2 U425 ( .A(n391), .B(n392), .S(n255), .Z(n390) );
  GTECH_NAND2 U426 ( .A(n393), .B(n296), .Z(n389) );
  GTECH_MUX2 U427 ( .A(n394), .B(n395), .S(n255), .Z(n393) );
  GTECH_NOT U428 ( .A(n391), .Z(n395) );
  GTECH_OAI22 U429 ( .A(n304), .B(n388), .C(n302), .D(n386), .Z(n391) );
  GTECH_NOT U430 ( .A(n392), .Z(n394) );
  GTECH_OAI22 U431 ( .A(n396), .B(n304), .C(n397), .D(n302), .Z(n392) );
  GTECH_NOT U432 ( .A(n386), .Z(n397) );
  GTECH_OAI21 U433 ( .A(n254), .B(n398), .C(n399), .Z(n386) );
  GTECH_OAI21 U434 ( .A(n35), .B(n400), .C(n401), .Z(n399) );
  GTECH_NOT U435 ( .A(n388), .Z(n396) );
  GTECH_OAI21 U436 ( .A(n35), .B(n254), .C(n402), .Z(n388) );
  GTECH_OAI21 U437 ( .A(n400), .B(n398), .C(n403), .Z(n402) );
  GTECH_NOT U438 ( .A(n35), .Z(n398) );
  GTECH_NOT U439 ( .A(n254), .Z(n400) );
  GTECH_AND2 U440 ( .A(n260), .B(n285), .Z(N109) );
  GTECH_MUX2 U441 ( .A(n404), .B(n405), .S(n35), .Z(n285) );
  GTECH_MUX2 U442 ( .A(n406), .B(n407), .S(n254), .Z(n405) );
  GTECH_NAND2 U443 ( .A(n408), .B(n296), .Z(n404) );
  GTECH_MUX2 U444 ( .A(n409), .B(n410), .S(n254), .Z(n408) );
  GTECH_NOT U445 ( .A(n406), .Z(n410) );
  GTECH_OAI22 U446 ( .A(n304), .B(n403), .C(n302), .D(n401), .Z(n406) );
  GTECH_NOT U447 ( .A(n407), .Z(n409) );
  GTECH_OAI22 U448 ( .A(n411), .B(n304), .C(n412), .D(n302), .Z(n407) );
  GTECH_NOT U449 ( .A(n401), .Z(n412) );
  GTECH_OAI21 U450 ( .A(n253), .B(n413), .C(n414), .Z(n401) );
  GTECH_OAI21 U451 ( .A(n36), .B(n415), .C(n416), .Z(n414) );
  GTECH_NOT U452 ( .A(n403), .Z(n411) );
  GTECH_OAI21 U453 ( .A(n36), .B(n253), .C(n417), .Z(n403) );
  GTECH_OAI21 U454 ( .A(n415), .B(n413), .C(n418), .Z(n417) );
  GTECH_NOT U455 ( .A(n36), .Z(n413) );
  GTECH_NOT U456 ( .A(n253), .Z(n415) );
  GTECH_AND2 U457 ( .A(n260), .B(n286), .Z(N108) );
  GTECH_MUX2 U458 ( .A(n419), .B(n420), .S(n36), .Z(n286) );
  GTECH_MUX2 U459 ( .A(n421), .B(n422), .S(n253), .Z(n420) );
  GTECH_NAND2 U460 ( .A(n423), .B(n296), .Z(n419) );
  GTECH_MUX2 U461 ( .A(n424), .B(n425), .S(n253), .Z(n423) );
  GTECH_NOT U462 ( .A(n421), .Z(n425) );
  GTECH_OAI22 U463 ( .A(n304), .B(n418), .C(n302), .D(n416), .Z(n421) );
  GTECH_NOT U464 ( .A(n422), .Z(n424) );
  GTECH_OAI22 U465 ( .A(n426), .B(n304), .C(n427), .D(n302), .Z(n422) );
  GTECH_NOT U466 ( .A(n416), .Z(n427) );
  GTECH_OAI21 U467 ( .A(n252), .B(n428), .C(n429), .Z(n416) );
  GTECH_OAI21 U468 ( .A(n37), .B(n430), .C(n431), .Z(n429) );
  GTECH_NOT U469 ( .A(n418), .Z(n426) );
  GTECH_OAI21 U470 ( .A(n37), .B(n252), .C(n432), .Z(n418) );
  GTECH_OAI21 U471 ( .A(n430), .B(n428), .C(n433), .Z(n432) );
  GTECH_NOT U472 ( .A(n37), .Z(n428) );
  GTECH_NOT U473 ( .A(n252), .Z(n430) );
  GTECH_AND2 U474 ( .A(n260), .B(n287), .Z(N107) );
  GTECH_MUX2 U475 ( .A(n434), .B(n435), .S(n37), .Z(n287) );
  GTECH_MUX2 U476 ( .A(n436), .B(n437), .S(n252), .Z(n435) );
  GTECH_NAND2 U477 ( .A(n438), .B(n296), .Z(n434) );
  GTECH_MUX2 U478 ( .A(n439), .B(n440), .S(n252), .Z(n438) );
  GTECH_NOT U479 ( .A(n436), .Z(n440) );
  GTECH_OAI22 U480 ( .A(n304), .B(n433), .C(n302), .D(n431), .Z(n436) );
  GTECH_NOT U481 ( .A(n437), .Z(n439) );
  GTECH_OAI22 U482 ( .A(n441), .B(n304), .C(n442), .D(n302), .Z(n437) );
  GTECH_NOT U483 ( .A(n431), .Z(n442) );
  GTECH_OAI21 U484 ( .A(n251), .B(n443), .C(n444), .Z(n431) );
  GTECH_OAI21 U485 ( .A(n38), .B(n445), .C(n446), .Z(n444) );
  GTECH_NOT U486 ( .A(n433), .Z(n441) );
  GTECH_OAI21 U487 ( .A(n38), .B(n251), .C(n447), .Z(n433) );
  GTECH_OAI21 U488 ( .A(n445), .B(n443), .C(n448), .Z(n447) );
  GTECH_NOT U489 ( .A(n38), .Z(n443) );
  GTECH_NOT U490 ( .A(n251), .Z(n445) );
  GTECH_AND2 U491 ( .A(n260), .B(n288), .Z(N106) );
  GTECH_MUX2 U492 ( .A(n449), .B(n450), .S(n38), .Z(n288) );
  GTECH_MUX2 U493 ( .A(n451), .B(n452), .S(n251), .Z(n450) );
  GTECH_NAND2 U494 ( .A(n453), .B(n296), .Z(n449) );
  GTECH_MUX2 U495 ( .A(n454), .B(n455), .S(n251), .Z(n453) );
  GTECH_NOT U496 ( .A(n451), .Z(n455) );
  GTECH_OAI22 U497 ( .A(n304), .B(n448), .C(n302), .D(n446), .Z(n451) );
  GTECH_NOT U498 ( .A(n452), .Z(n454) );
  GTECH_OAI22 U499 ( .A(n456), .B(n304), .C(n457), .D(n302), .Z(n452) );
  GTECH_NOT U500 ( .A(n446), .Z(n457) );
  GTECH_OAI21 U501 ( .A(n250), .B(n458), .C(n459), .Z(n446) );
  GTECH_OAI21 U502 ( .A(n39), .B(n460), .C(n461), .Z(n459) );
  GTECH_NOT U503 ( .A(n448), .Z(n456) );
  GTECH_OAI21 U504 ( .A(n39), .B(n250), .C(n462), .Z(n448) );
  GTECH_OAI21 U505 ( .A(n460), .B(n458), .C(n463), .Z(n462) );
  GTECH_NOT U506 ( .A(n39), .Z(n458) );
  GTECH_NOT U507 ( .A(n250), .Z(n460) );
  GTECH_AND2 U508 ( .A(n260), .B(n289), .Z(N105) );
  GTECH_MUX2 U509 ( .A(n464), .B(n465), .S(n39), .Z(n289) );
  GTECH_MUX2 U510 ( .A(n466), .B(n467), .S(n250), .Z(n465) );
  GTECH_NAND2 U511 ( .A(n468), .B(n296), .Z(n464) );
  GTECH_MUX2 U512 ( .A(n469), .B(n470), .S(n250), .Z(n468) );
  GTECH_NOT U513 ( .A(n466), .Z(n470) );
  GTECH_OAI22 U514 ( .A(n304), .B(n463), .C(n302), .D(n461), .Z(n466) );
  GTECH_NOT U515 ( .A(n467), .Z(n469) );
  GTECH_OAI22 U516 ( .A(n471), .B(n304), .C(n472), .D(n302), .Z(n467) );
  GTECH_NOT U517 ( .A(n461), .Z(n472) );
  GTECH_OAI21 U518 ( .A(n249), .B(n473), .C(n474), .Z(n461) );
  GTECH_OAI21 U519 ( .A(n40), .B(n475), .C(n476), .Z(n474) );
  GTECH_NOT U520 ( .A(n463), .Z(n471) );
  GTECH_OAI21 U521 ( .A(n40), .B(n249), .C(n477), .Z(n463) );
  GTECH_OAI21 U522 ( .A(n475), .B(n473), .C(n478), .Z(n477) );
  GTECH_NOT U523 ( .A(n40), .Z(n473) );
  GTECH_NOT U524 ( .A(n249), .Z(n475) );
  GTECH_AND2 U525 ( .A(n260), .B(n290), .Z(N104) );
  GTECH_MUX2 U526 ( .A(n479), .B(n480), .S(n40), .Z(n290) );
  GTECH_MUX2 U527 ( .A(n481), .B(n482), .S(n249), .Z(n480) );
  GTECH_NAND2 U528 ( .A(n483), .B(n296), .Z(n479) );
  GTECH_MUX2 U529 ( .A(n484), .B(n485), .S(n249), .Z(n483) );
  GTECH_NOT U530 ( .A(n481), .Z(n485) );
  GTECH_OAI22 U531 ( .A(n304), .B(n478), .C(n302), .D(n476), .Z(n481) );
  GTECH_NOT U532 ( .A(n482), .Z(n484) );
  GTECH_OAI22 U533 ( .A(n486), .B(n304), .C(n487), .D(n302), .Z(n482) );
  GTECH_NOT U534 ( .A(n476), .Z(n487) );
  GTECH_OAI21 U535 ( .A(n248), .B(n488), .C(n489), .Z(n476) );
  GTECH_OAI21 U536 ( .A(n41), .B(n490), .C(n491), .Z(n489) );
  GTECH_NOT U537 ( .A(n478), .Z(n486) );
  GTECH_OAI21 U538 ( .A(n41), .B(n248), .C(n492), .Z(n478) );
  GTECH_OAI21 U539 ( .A(n490), .B(n488), .C(n493), .Z(n492) );
  GTECH_NOT U540 ( .A(n41), .Z(n488) );
  GTECH_NOT U541 ( .A(n248), .Z(n490) );
  GTECH_AND2 U542 ( .A(n260), .B(n291), .Z(N103) );
  GTECH_MUX2 U543 ( .A(n494), .B(n495), .S(n41), .Z(n291) );
  GTECH_MUX2 U544 ( .A(n496), .B(n497), .S(n248), .Z(n495) );
  GTECH_NAND2 U545 ( .A(n498), .B(n296), .Z(n494) );
  GTECH_MUX2 U546 ( .A(n499), .B(n500), .S(n248), .Z(n498) );
  GTECH_NOT U547 ( .A(n496), .Z(n500) );
  GTECH_OAI22 U548 ( .A(n304), .B(n493), .C(n302), .D(n491), .Z(n496) );
  GTECH_NOT U549 ( .A(n497), .Z(n499) );
  GTECH_OAI22 U550 ( .A(n501), .B(n304), .C(n502), .D(n302), .Z(n497) );
  GTECH_NOT U551 ( .A(n491), .Z(n502) );
  GTECH_OAI21 U552 ( .A(n247), .B(n503), .C(n504), .Z(n491) );
  GTECH_OAI21 U553 ( .A(n42), .B(n505), .C(n506), .Z(n504) );
  GTECH_NOT U554 ( .A(n493), .Z(n501) );
  GTECH_OAI21 U555 ( .A(n42), .B(n247), .C(n507), .Z(n493) );
  GTECH_OAI21 U556 ( .A(n505), .B(n503), .C(n508), .Z(n507) );
  GTECH_NOT U557 ( .A(n42), .Z(n503) );
  GTECH_NOT U558 ( .A(n247), .Z(n505) );
  GTECH_AND2 U559 ( .A(n260), .B(n293), .Z(N102) );
  GTECH_MUX2 U560 ( .A(n509), .B(n510), .S(n42), .Z(n293) );
  GTECH_MUX2 U561 ( .A(n511), .B(n512), .S(n247), .Z(n510) );
  GTECH_NAND2 U562 ( .A(n513), .B(n296), .Z(n509) );
  GTECH_MUX2 U563 ( .A(n514), .B(n515), .S(n247), .Z(n513) );
  GTECH_NOT U564 ( .A(n511), .Z(n515) );
  GTECH_OAI22 U565 ( .A(n304), .B(n508), .C(n302), .D(n506), .Z(n511) );
  GTECH_NOT U566 ( .A(n512), .Z(n514) );
  GTECH_OAI22 U567 ( .A(n516), .B(n304), .C(n517), .D(n302), .Z(n512) );
  GTECH_NOT U568 ( .A(n506), .Z(n517) );
  GTECH_OAI21 U569 ( .A(n246), .B(n518), .C(n519), .Z(n506) );
  GTECH_OAI21 U570 ( .A(n43), .B(n520), .C(n521), .Z(n519) );
  GTECH_NOT U571 ( .A(n508), .Z(n516) );
  GTECH_OAI21 U572 ( .A(n43), .B(n246), .C(n522), .Z(n508) );
  GTECH_OAI21 U573 ( .A(n520), .B(n518), .C(n523), .Z(n522) );
  GTECH_NOT U574 ( .A(n43), .Z(n518) );
  GTECH_NOT U575 ( .A(n246), .Z(n520) );
  GTECH_AND2 U576 ( .A(n260), .B(n294), .Z(N101) );
  GTECH_MUX2 U577 ( .A(n524), .B(n525), .S(n43), .Z(n294) );
  GTECH_MUX2 U578 ( .A(n526), .B(n527), .S(n246), .Z(n525) );
  GTECH_NAND2 U579 ( .A(n528), .B(n296), .Z(n524) );
  GTECH_MUX2 U580 ( .A(n529), .B(n530), .S(n246), .Z(n528) );
  GTECH_NOT U581 ( .A(n526), .Z(n530) );
  GTECH_OAI22 U582 ( .A(n304), .B(n523), .C(n302), .D(n521), .Z(n526) );
  GTECH_NOT U583 ( .A(n527), .Z(n529) );
  GTECH_OAI22 U584 ( .A(n531), .B(n304), .C(n532), .D(n302), .Z(n527) );
  GTECH_NOT U585 ( .A(n521), .Z(n532) );
  GTECH_OAI21 U586 ( .A(n245), .B(n533), .C(n534), .Z(n521) );
  GTECH_OAI21 U587 ( .A(n29), .B(n535), .C(n536), .Z(n534) );
  GTECH_NOT U588 ( .A(n523), .Z(n531) );
  GTECH_OAI21 U589 ( .A(n29), .B(n245), .C(n537), .Z(n523) );
  GTECH_OAI21 U590 ( .A(n535), .B(n533), .C(n538), .Z(n537) );
  GTECH_NOT U591 ( .A(n29), .Z(n533) );
  GTECH_NOT U592 ( .A(n245), .Z(n535) );
  GTECH_AND2 U593 ( .A(n260), .B(n295), .Z(N100) );
  GTECH_MUX2 U594 ( .A(n539), .B(n540), .S(n29), .Z(n295) );
  GTECH_MUX2 U595 ( .A(n541), .B(n542), .S(n245), .Z(n540) );
  GTECH_NAND2 U596 ( .A(n543), .B(n296), .Z(n539) );
  GTECH_NAND2 U597 ( .A(n304), .B(n302), .Z(n296) );
  GTECH_MUX2 U598 ( .A(n544), .B(n545), .S(n245), .Z(n543) );
  GTECH_NOT U599 ( .A(n541), .Z(n545) );
  GTECH_OAI22 U600 ( .A(n304), .B(n538), .C(n302), .D(n536), .Z(n541) );
  GTECH_NOT U601 ( .A(n542), .Z(n544) );
  GTECH_OAI22 U602 ( .A(n546), .B(n304), .C(n547), .D(n302), .Z(n542) );
  GTECH_NAND2 U603 ( .A(n10), .B(n265), .Z(n302) );
  GTECH_NOT U604 ( .A(n28), .Z(n265) );
  GTECH_NOT U605 ( .A(n536), .Z(n547) );
  GTECH_OAI21 U606 ( .A(n244), .B(n548), .C(n549), .Z(n536) );
  GTECH_OAI21 U607 ( .A(n11), .B(n550), .C(n301), .Z(n549) );
  GTECH_NOT U608 ( .A(n305), .Z(n301) );
  GTECH_NAND2 U609 ( .A(n12), .B(n309), .Z(n305) );
  GTECH_NAND2 U610 ( .A(n28), .B(n551), .Z(n304) );
  GTECH_NOT U611 ( .A(n10), .Z(n551) );
  GTECH_NOT U612 ( .A(n538), .Z(n546) );
  GTECH_OAI21 U613 ( .A(n244), .B(n11), .C(n552), .Z(n538) );
  GTECH_OAI21 U614 ( .A(n550), .B(n548), .C(n303), .Z(n552) );
  GTECH_NOT U615 ( .A(n306), .Z(n303) );
  GTECH_NAND2 U616 ( .A(n553), .B(n309), .Z(n306) );
  GTECH_NOT U617 ( .A(n243), .Z(n309) );
  GTECH_NOT U618 ( .A(n12), .Z(n553) );
  GTECH_NOT U619 ( .A(n11), .Z(n548) );
  GTECH_NOT U620 ( .A(n244), .Z(n550) );
  GTECH_NOT U621 ( .A(n263), .Z(n260) );
  GTECH_OAI21 U622 ( .A(n268), .B(n269), .C(n270), .Z(n263) );
  GTECH_NOT U623 ( .A(n554), .Z(n270) );
  GTECH_NAND2 U624 ( .A(n277), .B(n555), .Z(n554) );
  GTECH_NOT U625 ( .A(Ld), .Z(n555) );
  GTECH_NOT U626 ( .A(Rst), .Z(n277) );
  GTECH_NOT U627 ( .A(n9), .Z(n269) );
  GTECH_NAND2 U628 ( .A(n8), .B(n272), .Z(n268) );
  GTECH_NOT U629 ( .A(n275), .Z(n272) );
  GTECH_NAND2 U630 ( .A(n7), .B(n274), .Z(n275) );
  GTECH_NOT U631 ( .A(n556), .Z(n274) );
  GTECH_NAND2 U632 ( .A(n6), .B(n242), .Z(n556) );
endmodule

