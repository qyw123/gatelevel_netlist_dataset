
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371;

  GTECH_MUX2 U134 ( .A(n273), .B(n274), .S(n275), .Z(sum[9]) );
  GTECH_XOR2 U135 ( .A(n276), .B(n277), .Z(n274) );
  GTECH_XOR2 U136 ( .A(n278), .B(n277), .Z(n273) );
  GTECH_OAI21 U137 ( .A(a[9]), .B(b[9]), .C(n279), .Z(n277) );
  GTECH_NAND2 U138 ( .A(n280), .B(n281), .Z(sum[8]) );
  GTECH_AO21 U139 ( .A(n276), .B(n282), .C(n275), .Z(n280) );
  GTECH_MUX2 U140 ( .A(n283), .B(n284), .S(n285), .Z(sum[7]) );
  GTECH_XOR2 U141 ( .A(n286), .B(n287), .Z(n284) );
  GTECH_OA21 U142 ( .A(n288), .B(n289), .C(n290), .Z(n287) );
  GTECH_XNOR2 U143 ( .A(n286), .B(n291), .Z(n283) );
  GTECH_XNOR2 U144 ( .A(a[7]), .B(b[7]), .Z(n286) );
  GTECH_MUX2 U145 ( .A(n292), .B(n293), .S(n285), .Z(sum[6]) );
  GTECH_XNOR2 U146 ( .A(n294), .B(n289), .Z(n293) );
  GTECH_OA21 U147 ( .A(n295), .B(n296), .C(n297), .Z(n289) );
  GTECH_XNOR2 U148 ( .A(n294), .B(n298), .Z(n292) );
  GTECH_AND_NOT U149 ( .A(n290), .B(n288), .Z(n294) );
  GTECH_XNOR2 U150 ( .A(n299), .B(n300), .Z(sum[5]) );
  GTECH_OA21 U151 ( .A(n301), .B(n285), .C(n296), .Z(n300) );
  GTECH_AND_NOT U152 ( .A(n297), .B(n295), .Z(n299) );
  GTECH_XNOR2 U153 ( .A(n302), .B(n285), .Z(sum[4]) );
  GTECH_MUX2 U154 ( .A(n303), .B(n304), .S(cin), .Z(sum[3]) );
  GTECH_XNOR2 U155 ( .A(n305), .B(n306), .Z(n304) );
  GTECH_XOR2 U156 ( .A(n305), .B(n307), .Z(n303) );
  GTECH_AOI21 U157 ( .A(n308), .B(n309), .C(n310), .Z(n307) );
  GTECH_XNOR2 U158 ( .A(a[3]), .B(b[3]), .Z(n305) );
  GTECH_MUX2 U159 ( .A(n311), .B(n312), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U160 ( .A(n313), .B(n314), .Z(n312) );
  GTECH_XOR2 U161 ( .A(n309), .B(n313), .Z(n311) );
  GTECH_AND_NOT U162 ( .A(n308), .B(n310), .Z(n313) );
  GTECH_OAI21 U163 ( .A(n315), .B(n316), .C(n317), .Z(n309) );
  GTECH_MUX2 U164 ( .A(n318), .B(n319), .S(n320), .Z(sum[1]) );
  GTECH_AND_NOT U165 ( .A(n317), .B(n315), .Z(n320) );
  GTECH_AO21 U166 ( .A(n321), .B(n316), .C(n322), .Z(n319) );
  GTECH_OAI21 U167 ( .A(n322), .B(n321), .C(n316), .Z(n318) );
  GTECH_NAND2 U168 ( .A(a[0]), .B(b[0]), .Z(n316) );
  GTECH_NOT U169 ( .A(cin), .Z(n321) );
  GTECH_MUX2 U170 ( .A(n323), .B(n324), .S(n325), .Z(sum[15]) );
  GTECH_XOR2 U171 ( .A(n326), .B(n327), .Z(n324) );
  GTECH_AOI21 U172 ( .A(n328), .B(n329), .C(n330), .Z(n327) );
  GTECH_XNOR2 U173 ( .A(n326), .B(n331), .Z(n323) );
  GTECH_XNOR2 U174 ( .A(a[15]), .B(b[15]), .Z(n326) );
  GTECH_MUX2 U175 ( .A(n332), .B(n333), .S(n325), .Z(sum[14]) );
  GTECH_XOR2 U176 ( .A(n334), .B(n329), .Z(n333) );
  GTECH_AOI21 U177 ( .A(n335), .B(n336), .C(n337), .Z(n329) );
  GTECH_XOR2 U178 ( .A(n334), .B(n338), .Z(n332) );
  GTECH_AND_NOT U179 ( .A(n328), .B(n330), .Z(n334) );
  GTECH_MUX2 U180 ( .A(n339), .B(n340), .S(n325), .Z(sum[13]) );
  GTECH_XNOR2 U181 ( .A(n341), .B(n342), .Z(n340) );
  GTECH_XOR2 U182 ( .A(n342), .B(n343), .Z(n339) );
  GTECH_OAI21 U183 ( .A(a[13]), .B(b[13]), .C(n335), .Z(n342) );
  GTECH_NAND2 U184 ( .A(n344), .B(n345), .Z(sum[12]) );
  GTECH_OAI21 U185 ( .A(n341), .B(n343), .C(n346), .Z(n344) );
  GTECH_MUX2 U186 ( .A(n347), .B(n348), .S(n275), .Z(sum[11]) );
  GTECH_XOR2 U187 ( .A(n349), .B(n350), .Z(n348) );
  GTECH_AOI21 U188 ( .A(n351), .B(n352), .C(n353), .Z(n350) );
  GTECH_XNOR2 U189 ( .A(n349), .B(n354), .Z(n347) );
  GTECH_XNOR2 U190 ( .A(a[11]), .B(b[11]), .Z(n349) );
  GTECH_MUX2 U191 ( .A(n355), .B(n356), .S(n275), .Z(sum[10]) );
  GTECH_XOR2 U192 ( .A(n357), .B(n352), .Z(n356) );
  GTECH_AOI21 U193 ( .A(n279), .B(n276), .C(n358), .Z(n352) );
  GTECH_XOR2 U194 ( .A(n357), .B(n359), .Z(n355) );
  GTECH_AND_NOT U195 ( .A(n351), .B(n353), .Z(n357) );
  GTECH_XNOR2 U196 ( .A(cin), .B(n360), .Z(sum[0]) );
  GTECH_OAI21 U197 ( .A(n325), .B(n361), .C(n345), .Z(cout) );
  GTECH_OR3 U198 ( .A(n341), .B(n343), .C(n346), .Z(n345) );
  GTECH_NOT U199 ( .A(n336), .Z(n341) );
  GTECH_NAND2 U200 ( .A(a[12]), .B(b[12]), .Z(n336) );
  GTECH_AOI21 U201 ( .A(n331), .B(a[15]), .C(n362), .Z(n361) );
  GTECH_OA21 U202 ( .A(a[15]), .B(n331), .C(b[15]), .Z(n362) );
  GTECH_AO21 U203 ( .A(n328), .B(n338), .C(n330), .Z(n331) );
  GTECH_AND2 U204 ( .A(a[14]), .B(b[14]), .Z(n330) );
  GTECH_AOI21 U205 ( .A(n335), .B(n343), .C(n337), .Z(n338) );
  GTECH_NOR2 U206 ( .A(b[13]), .B(a[13]), .Z(n337) );
  GTECH_NOR2 U207 ( .A(b[12]), .B(a[12]), .Z(n343) );
  GTECH_NAND2 U208 ( .A(a[13]), .B(b[13]), .Z(n335) );
  GTECH_OR2 U209 ( .A(a[14]), .B(b[14]), .Z(n328) );
  GTECH_NOT U210 ( .A(n346), .Z(n325) );
  GTECH_OAI21 U211 ( .A(n363), .B(n275), .C(n281), .Z(n346) );
  GTECH_NAND3 U212 ( .A(n282), .B(n276), .C(n275), .Z(n281) );
  GTECH_NAND2 U213 ( .A(b[8]), .B(a[8]), .Z(n276) );
  GTECH_NOT U214 ( .A(n278), .Z(n282) );
  GTECH_NOT U215 ( .A(n364), .Z(n275) );
  GTECH_MUX2 U216 ( .A(n365), .B(n302), .S(n285), .Z(n364) );
  GTECH_MUX2 U217 ( .A(n360), .B(n366), .S(cin), .Z(n285) );
  GTECH_AOI21 U218 ( .A(n306), .B(a[3]), .C(n367), .Z(n366) );
  GTECH_OA21 U219 ( .A(a[3]), .B(n306), .C(b[3]), .Z(n367) );
  GTECH_AO21 U220 ( .A(n314), .B(n308), .C(n310), .Z(n306) );
  GTECH_AND2 U221 ( .A(b[2]), .B(a[2]), .Z(n310) );
  GTECH_OR2 U222 ( .A(a[2]), .B(b[2]), .Z(n308) );
  GTECH_OAI21 U223 ( .A(n322), .B(n315), .C(n317), .Z(n314) );
  GTECH_NAND2 U224 ( .A(b[1]), .B(a[1]), .Z(n317) );
  GTECH_NOR2 U225 ( .A(b[1]), .B(a[1]), .Z(n315) );
  GTECH_AND_NOT U226 ( .A(n368), .B(a[0]), .Z(n322) );
  GTECH_XNOR2 U227 ( .A(n369), .B(n368), .Z(n360) );
  GTECH_NOT U228 ( .A(b[0]), .Z(n368) );
  GTECH_NOT U229 ( .A(a[0]), .Z(n369) );
  GTECH_AND_NOT U230 ( .A(n296), .B(n301), .Z(n302) );
  GTECH_NAND2 U231 ( .A(b[4]), .B(a[4]), .Z(n296) );
  GTECH_OA21 U232 ( .A(a[7]), .B(n291), .C(n370), .Z(n365) );
  GTECH_AO21 U233 ( .A(n291), .B(a[7]), .C(b[7]), .Z(n370) );
  GTECH_OAI21 U234 ( .A(n298), .B(n288), .C(n290), .Z(n291) );
  GTECH_NAND2 U235 ( .A(b[6]), .B(a[6]), .Z(n290) );
  GTECH_NOR2 U236 ( .A(a[6]), .B(b[6]), .Z(n288) );
  GTECH_OA21 U237 ( .A(n301), .B(n295), .C(n297), .Z(n298) );
  GTECH_NAND2 U238 ( .A(b[5]), .B(a[5]), .Z(n297) );
  GTECH_NOR2 U239 ( .A(b[5]), .B(a[5]), .Z(n295) );
  GTECH_NOR2 U240 ( .A(a[4]), .B(b[4]), .Z(n301) );
  GTECH_AOI21 U241 ( .A(n354), .B(a[11]), .C(n371), .Z(n363) );
  GTECH_OA21 U242 ( .A(a[11]), .B(n354), .C(b[11]), .Z(n371) );
  GTECH_AO21 U243 ( .A(n351), .B(n359), .C(n353), .Z(n354) );
  GTECH_AND2 U244 ( .A(a[10]), .B(b[10]), .Z(n353) );
  GTECH_AOI21 U245 ( .A(n279), .B(n278), .C(n358), .Z(n359) );
  GTECH_NOR2 U246 ( .A(b[9]), .B(a[9]), .Z(n358) );
  GTECH_NOR2 U247 ( .A(a[8]), .B(b[8]), .Z(n278) );
  GTECH_NAND2 U248 ( .A(b[9]), .B(a[9]), .Z(n279) );
  GTECH_OR2 U249 ( .A(a[10]), .B(b[10]), .Z(n351) );
endmodule

