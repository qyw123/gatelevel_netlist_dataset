
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382;

  GTECH_MUX2 U140 ( .A(n279), .B(n280), .S(n281), .Z(sum[9]) );
  GTECH_XNOR2 U141 ( .A(n282), .B(n283), .Z(n280) );
  GTECH_XNOR2 U142 ( .A(n282), .B(n284), .Z(n279) );
  GTECH_AOI21 U143 ( .A(a[9]), .B(b[9]), .C(n285), .Z(n282) );
  GTECH_NAND2 U144 ( .A(n286), .B(n287), .Z(sum[8]) );
  GTECH_OAI21 U145 ( .A(n288), .B(n283), .C(n281), .Z(n286) );
  GTECH_MUX2 U146 ( .A(n289), .B(n290), .S(n291), .Z(sum[7]) );
  GTECH_XOR2 U147 ( .A(n292), .B(n293), .Z(n290) );
  GTECH_XNOR2 U148 ( .A(n292), .B(n294), .Z(n289) );
  GTECH_OA21 U149 ( .A(n295), .B(n296), .C(n297), .Z(n294) );
  GTECH_XOR2 U150 ( .A(a[7]), .B(b[7]), .Z(n292) );
  GTECH_MUX2 U151 ( .A(n298), .B(n299), .S(n300), .Z(sum[6]) );
  GTECH_OA21 U152 ( .A(n301), .B(n302), .C(n296), .Z(n300) );
  GTECH_OAI21 U153 ( .A(n303), .B(n304), .C(n305), .Z(n296) );
  GTECH_XOR2 U154 ( .A(b[6]), .B(a[6]), .Z(n299) );
  GTECH_OR_NOT U155 ( .A(n295), .B(n297), .Z(n298) );
  GTECH_XOR2 U156 ( .A(n306), .B(n307), .Z(sum[5]) );
  GTECH_OA21 U157 ( .A(n303), .B(n291), .C(n308), .Z(n307) );
  GTECH_AND_NOT U158 ( .A(n305), .B(n304), .Z(n306) );
  GTECH_XNOR2 U159 ( .A(n309), .B(n291), .Z(sum[4]) );
  GTECH_MUX2 U160 ( .A(n310), .B(n311), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U161 ( .A(n312), .B(n313), .Z(n311) );
  GTECH_XNOR2 U162 ( .A(n312), .B(n314), .Z(n310) );
  GTECH_AND2 U163 ( .A(n315), .B(n316), .Z(n314) );
  GTECH_OAI21 U164 ( .A(b[2]), .B(a[2]), .C(n317), .Z(n315) );
  GTECH_XOR2 U165 ( .A(a[3]), .B(b[3]), .Z(n312) );
  GTECH_MUX2 U166 ( .A(n318), .B(n319), .S(n320), .Z(sum[2]) );
  GTECH_NOT U167 ( .A(cin), .Z(n320) );
  GTECH_MUX2 U168 ( .A(n321), .B(n322), .S(n317), .Z(n319) );
  GTECH_OA21 U169 ( .A(n323), .B(n324), .C(n325), .Z(n317) );
  GTECH_MUX2 U170 ( .A(n321), .B(n322), .S(n326), .Z(n318) );
  GTECH_OAI21 U171 ( .A(b[2]), .B(a[2]), .C(n316), .Z(n322) );
  GTECH_XOR2 U172 ( .A(a[2]), .B(b[2]), .Z(n321) );
  GTECH_MUX2 U173 ( .A(n327), .B(n328), .S(n329), .Z(sum[1]) );
  GTECH_AND_NOT U174 ( .A(n325), .B(n324), .Z(n329) );
  GTECH_OAI21 U175 ( .A(cin), .B(n323), .C(n330), .Z(n328) );
  GTECH_AO21 U176 ( .A(n330), .B(cin), .C(n323), .Z(n327) );
  GTECH_AND2 U177 ( .A(b[0]), .B(a[0]), .Z(n323) );
  GTECH_MUX2 U178 ( .A(n331), .B(n332), .S(n333), .Z(sum[15]) );
  GTECH_XOR2 U179 ( .A(n334), .B(n335), .Z(n332) );
  GTECH_AND2 U180 ( .A(n336), .B(n337), .Z(n335) );
  GTECH_OAI21 U181 ( .A(b[14]), .B(a[14]), .C(n338), .Z(n336) );
  GTECH_XNOR2 U182 ( .A(n334), .B(n339), .Z(n331) );
  GTECH_XNOR2 U183 ( .A(a[15]), .B(b[15]), .Z(n334) );
  GTECH_OAI21 U184 ( .A(n340), .B(n337), .C(n341), .Z(sum[14]) );
  GTECH_MUX2 U185 ( .A(n342), .B(n343), .S(b[14]), .Z(n341) );
  GTECH_OR_NOT U186 ( .A(a[14]), .B(n340), .Z(n343) );
  GTECH_XOR2 U187 ( .A(a[14]), .B(n340), .Z(n342) );
  GTECH_AOI21 U188 ( .A(n344), .B(n345), .C(n338), .Z(n340) );
  GTECH_OAI2N2 U189 ( .A(n346), .B(n347), .C(a[13]), .D(b[13]), .Z(n338) );
  GTECH_MUX2 U190 ( .A(n348), .B(n349), .S(n333), .Z(sum[13]) );
  GTECH_XNOR2 U191 ( .A(n350), .B(n347), .Z(n349) );
  GTECH_XNOR2 U192 ( .A(n351), .B(n350), .Z(n348) );
  GTECH_AOI21 U193 ( .A(a[13]), .B(b[13]), .C(n346), .Z(n350) );
  GTECH_NAND2 U194 ( .A(n352), .B(n353), .Z(sum[12]) );
  GTECH_AO21 U195 ( .A(n347), .B(n354), .C(n333), .Z(n352) );
  GTECH_NOT U196 ( .A(n351), .Z(n354) );
  GTECH_NOT U197 ( .A(n355), .Z(n347) );
  GTECH_MUX2 U198 ( .A(n356), .B(n357), .S(n281), .Z(sum[11]) );
  GTECH_XOR2 U199 ( .A(n358), .B(n359), .Z(n357) );
  GTECH_XNOR2 U200 ( .A(n358), .B(n360), .Z(n356) );
  GTECH_AND2 U201 ( .A(n361), .B(n362), .Z(n360) );
  GTECH_OAI21 U202 ( .A(b[10]), .B(a[10]), .C(n363), .Z(n361) );
  GTECH_XOR2 U203 ( .A(a[11]), .B(b[11]), .Z(n358) );
  GTECH_OAI21 U204 ( .A(n364), .B(n362), .C(n365), .Z(sum[10]) );
  GTECH_MUX2 U205 ( .A(n366), .B(n367), .S(b[10]), .Z(n365) );
  GTECH_OR_NOT U206 ( .A(a[10]), .B(n364), .Z(n367) );
  GTECH_XOR2 U207 ( .A(a[10]), .B(n364), .Z(n366) );
  GTECH_AOI21 U208 ( .A(n368), .B(n281), .C(n363), .Z(n364) );
  GTECH_OAI2N2 U209 ( .A(n285), .B(n284), .C(a[9]), .D(b[9]), .Z(n363) );
  GTECH_NOT U210 ( .A(n288), .Z(n284) );
  GTECH_XNOR2 U211 ( .A(cin), .B(n369), .Z(sum[0]) );
  GTECH_OAI21 U212 ( .A(n333), .B(n370), .C(n353), .Z(cout) );
  GTECH_OR3 U213 ( .A(n355), .B(n351), .C(n344), .Z(n353) );
  GTECH_AND2 U214 ( .A(a[12]), .B(b[12]), .Z(n355) );
  GTECH_AOI21 U215 ( .A(n339), .B(a[15]), .C(n371), .Z(n370) );
  GTECH_OA21 U216 ( .A(a[15]), .B(n339), .C(b[15]), .Z(n371) );
  GTECH_NAND2 U217 ( .A(n372), .B(n337), .Z(n339) );
  GTECH_NAND2 U218 ( .A(a[14]), .B(b[14]), .Z(n337) );
  GTECH_OAI21 U219 ( .A(a[14]), .B(b[14]), .C(n345), .Z(n372) );
  GTECH_OAI2N2 U220 ( .A(n351), .B(n346), .C(a[13]), .D(b[13]), .Z(n345) );
  GTECH_NOR2 U221 ( .A(b[13]), .B(a[13]), .Z(n346) );
  GTECH_NOR2 U222 ( .A(b[12]), .B(a[12]), .Z(n351) );
  GTECH_NOT U223 ( .A(n344), .Z(n333) );
  GTECH_OAI21 U224 ( .A(n373), .B(n374), .C(n287), .Z(n344) );
  GTECH_OR3 U225 ( .A(n288), .B(n283), .C(n281), .Z(n287) );
  GTECH_NOT U226 ( .A(n374), .Z(n281) );
  GTECH_AND2 U227 ( .A(b[8]), .B(a[8]), .Z(n288) );
  GTECH_MUX2 U228 ( .A(n309), .B(n375), .S(n291), .Z(n374) );
  GTECH_NOT U229 ( .A(n301), .Z(n291) );
  GTECH_MUX2 U230 ( .A(n369), .B(n376), .S(cin), .Z(n301) );
  GTECH_AOI21 U231 ( .A(n313), .B(a[3]), .C(n377), .Z(n376) );
  GTECH_OA21 U232 ( .A(a[3]), .B(n313), .C(b[3]), .Z(n377) );
  GTECH_NAND2 U233 ( .A(n316), .B(n378), .Z(n313) );
  GTECH_OAI21 U234 ( .A(a[2]), .B(b[2]), .C(n326), .Z(n378) );
  GTECH_OA21 U235 ( .A(n324), .B(n330), .C(n325), .Z(n326) );
  GTECH_OR2 U236 ( .A(b[1]), .B(a[1]), .Z(n325) );
  GTECH_OR2 U237 ( .A(a[0]), .B(b[0]), .Z(n330) );
  GTECH_AND2 U238 ( .A(a[1]), .B(b[1]), .Z(n324) );
  GTECH_NAND2 U239 ( .A(b[2]), .B(a[2]), .Z(n316) );
  GTECH_XNOR2 U240 ( .A(a[0]), .B(b[0]), .Z(n369) );
  GTECH_AOI21 U241 ( .A(n293), .B(a[7]), .C(n379), .Z(n375) );
  GTECH_OA21 U242 ( .A(a[7]), .B(n293), .C(b[7]), .Z(n379) );
  GTECH_OAI21 U243 ( .A(n295), .B(n302), .C(n297), .Z(n293) );
  GTECH_OR_NOT U244 ( .A(n380), .B(b[6]), .Z(n297) );
  GTECH_NOT U245 ( .A(a[6]), .Z(n380) );
  GTECH_OAI21 U246 ( .A(n304), .B(n308), .C(n305), .Z(n302) );
  GTECH_OR2 U247 ( .A(a[5]), .B(b[5]), .Z(n305) );
  GTECH_AND2 U248 ( .A(b[5]), .B(a[5]), .Z(n304) );
  GTECH_NOR2 U249 ( .A(a[6]), .B(b[6]), .Z(n295) );
  GTECH_OR_NOT U250 ( .A(n303), .B(n308), .Z(n309) );
  GTECH_OR2 U251 ( .A(b[4]), .B(a[4]), .Z(n308) );
  GTECH_AND2 U252 ( .A(b[4]), .B(a[4]), .Z(n303) );
  GTECH_AOI21 U253 ( .A(n359), .B(a[11]), .C(n381), .Z(n373) );
  GTECH_OA21 U254 ( .A(a[11]), .B(n359), .C(b[11]), .Z(n381) );
  GTECH_NAND2 U255 ( .A(n382), .B(n362), .Z(n359) );
  GTECH_NAND2 U256 ( .A(a[10]), .B(b[10]), .Z(n362) );
  GTECH_OAI21 U257 ( .A(a[10]), .B(b[10]), .C(n368), .Z(n382) );
  GTECH_OAI2N2 U258 ( .A(n283), .B(n285), .C(a[9]), .D(b[9]), .Z(n368) );
  GTECH_NOR2 U259 ( .A(a[9]), .B(b[9]), .Z(n285) );
  GTECH_NOR2 U260 ( .A(a[8]), .B(b[8]), .Z(n283) );
endmodule

