
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393;

  GTECH_MUX2 U139 ( .A(n278), .B(n279), .S(n280), .Z(sum[9]) );
  GTECH_XOR2 U140 ( .A(n281), .B(n282), .Z(n279) );
  GTECH_NOT U141 ( .A(n283), .Z(n282) );
  GTECH_XOR2 U142 ( .A(n281), .B(n284), .Z(n278) );
  GTECH_AOI21 U143 ( .A(a[9]), .B(b[9]), .C(n285), .Z(n281) );
  GTECH_XOR2 U144 ( .A(n280), .B(n286), .Z(sum[8]) );
  GTECH_MUX2 U145 ( .A(n287), .B(n288), .S(n289), .Z(sum[7]) );
  GTECH_XOR2 U146 ( .A(n290), .B(n291), .Z(n288) );
  GTECH_XNOR2 U147 ( .A(n290), .B(n292), .Z(n287) );
  GTECH_OA21 U148 ( .A(n293), .B(n294), .C(n295), .Z(n292) );
  GTECH_XOR2 U149 ( .A(a[7]), .B(b[7]), .Z(n290) );
  GTECH_OAI21 U150 ( .A(n296), .B(n295), .C(n297), .Z(sum[6]) );
  GTECH_MUX2 U151 ( .A(n298), .B(n299), .S(b[6]), .Z(n297) );
  GTECH_OR_NOT U152 ( .A(a[6]), .B(n296), .Z(n299) );
  GTECH_XNOR2 U153 ( .A(n300), .B(n296), .Z(n298) );
  GTECH_OA21 U154 ( .A(n301), .B(n302), .C(n294), .Z(n296) );
  GTECH_AOI21 U155 ( .A(n303), .B(n304), .C(n305), .Z(n294) );
  GTECH_MUX2 U156 ( .A(n306), .B(n307), .S(n308), .Z(sum[5]) );
  GTECH_AND_NOT U157 ( .A(n303), .B(n305), .Z(n308) );
  GTECH_OAI22 U158 ( .A(n304), .B(n289), .C(b[4]), .D(a[4]), .Z(n307) );
  GTECH_ADD_AB U159 ( .A(b[4]), .B(a[4]), .COUT(n304) );
  GTECH_AO21 U160 ( .A(n289), .B(a[4]), .C(n309), .Z(n306) );
  GTECH_NOT U161 ( .A(n310), .Z(n309) );
  GTECH_OAI21 U162 ( .A(a[4]), .B(n289), .C(b[4]), .Z(n310) );
  GTECH_XNOR2 U163 ( .A(n311), .B(n302), .Z(sum[4]) );
  GTECH_NOT U164 ( .A(n289), .Z(n302) );
  GTECH_MUX2 U165 ( .A(n312), .B(n313), .S(n314), .Z(sum[3]) );
  GTECH_XNOR2 U166 ( .A(n315), .B(n316), .Z(n313) );
  GTECH_OA21 U167 ( .A(n317), .B(n318), .C(n319), .Z(n316) );
  GTECH_XOR2 U168 ( .A(n315), .B(n320), .Z(n312) );
  GTECH_XOR2 U169 ( .A(a[3]), .B(b[3]), .Z(n315) );
  GTECH_MUX2 U170 ( .A(n321), .B(n322), .S(cin), .Z(sum[2]) );
  GTECH_MUX2 U171 ( .A(n323), .B(n324), .S(n325), .Z(n322) );
  GTECH_MUX2 U172 ( .A(n323), .B(n324), .S(n318), .Z(n321) );
  GTECH_AOI21 U173 ( .A(n326), .B(n327), .C(n328), .Z(n318) );
  GTECH_XOR2 U174 ( .A(n329), .B(n330), .Z(n324) );
  GTECH_OAI21 U175 ( .A(b[2]), .B(a[2]), .C(n319), .Z(n323) );
  GTECH_MUX2 U176 ( .A(n331), .B(n332), .S(n333), .Z(sum[1]) );
  GTECH_AND_NOT U177 ( .A(n326), .B(n328), .Z(n333) );
  GTECH_OAI21 U178 ( .A(cin), .B(n327), .C(n334), .Z(n332) );
  GTECH_AO21 U179 ( .A(n334), .B(cin), .C(n327), .Z(n331) );
  GTECH_MUX2 U180 ( .A(n335), .B(n336), .S(n337), .Z(sum[15]) );
  GTECH_XOR2 U181 ( .A(n338), .B(n339), .Z(n336) );
  GTECH_OA21 U182 ( .A(n340), .B(n341), .C(n342), .Z(n339) );
  GTECH_XOR2 U183 ( .A(n338), .B(n343), .Z(n335) );
  GTECH_NOT U184 ( .A(n344), .Z(n343) );
  GTECH_XNOR2 U185 ( .A(a[15]), .B(b[15]), .Z(n338) );
  GTECH_OAI21 U186 ( .A(n345), .B(n342), .C(n346), .Z(sum[14]) );
  GTECH_MUX2 U187 ( .A(n347), .B(n348), .S(n349), .Z(n346) );
  GTECH_XOR2 U188 ( .A(a[14]), .B(n345), .Z(n348) );
  GTECH_OR_NOT U189 ( .A(a[14]), .B(n345), .Z(n347) );
  GTECH_OA21 U190 ( .A(n337), .B(n350), .C(n341), .Z(n345) );
  GTECH_OAI21 U191 ( .A(n351), .B(n352), .C(n353), .Z(n341) );
  GTECH_MUX2 U192 ( .A(n354), .B(n355), .S(n337), .Z(sum[13]) );
  GTECH_XOR2 U193 ( .A(n351), .B(n356), .Z(n355) );
  GTECH_XOR2 U194 ( .A(n357), .B(n356), .Z(n354) );
  GTECH_OA21 U195 ( .A(a[13]), .B(b[13]), .C(n358), .Z(n356) );
  GTECH_NOT U196 ( .A(n352), .Z(n358) );
  GTECH_XOR2 U197 ( .A(n359), .B(n337), .Z(sum[12]) );
  GTECH_MUX2 U198 ( .A(n360), .B(n361), .S(n280), .Z(sum[11]) );
  GTECH_XOR2 U199 ( .A(n362), .B(n363), .Z(n361) );
  GTECH_XNOR2 U200 ( .A(n362), .B(n364), .Z(n360) );
  GTECH_OA21 U201 ( .A(n365), .B(n366), .C(n367), .Z(n364) );
  GTECH_XOR2 U202 ( .A(a[11]), .B(b[11]), .Z(n362) );
  GTECH_OAI21 U203 ( .A(n368), .B(n367), .C(n369), .Z(sum[10]) );
  GTECH_MUX2 U204 ( .A(n370), .B(n371), .S(b[10]), .Z(n369) );
  GTECH_OR_NOT U205 ( .A(a[10]), .B(n368), .Z(n371) );
  GTECH_XOR2 U206 ( .A(a[10]), .B(n368), .Z(n370) );
  GTECH_OA21 U207 ( .A(n372), .B(n373), .C(n366), .Z(n368) );
  GTECH_AOI22 U208 ( .A(a[9]), .B(b[9]), .C(n374), .D(n284), .Z(n366) );
  GTECH_NOT U209 ( .A(n280), .Z(n373) );
  GTECH_XNOR2 U210 ( .A(n314), .B(n375), .Z(sum[0]) );
  GTECH_NOT U211 ( .A(n376), .Z(cout) );
  GTECH_MUX2 U212 ( .A(n377), .B(n359), .S(n337), .Z(n376) );
  GTECH_MUX2 U213 ( .A(n378), .B(n379), .S(n280), .Z(n337) );
  GTECH_MUX2 U214 ( .A(n311), .B(n380), .S(n289), .Z(n280) );
  GTECH_MUX2 U215 ( .A(n381), .B(n375), .S(n314), .Z(n289) );
  GTECH_NOT U216 ( .A(cin), .Z(n314) );
  GTECH_AND_NOT U217 ( .A(n334), .B(n327), .Z(n375) );
  GTECH_ADD_AB U218 ( .A(a[0]), .B(b[0]), .COUT(n327) );
  GTECH_OA21 U219 ( .A(a[3]), .B(n320), .C(n382), .Z(n381) );
  GTECH_AO21 U220 ( .A(n320), .B(a[3]), .C(b[3]), .Z(n382) );
  GTECH_OAI21 U221 ( .A(n325), .B(n317), .C(n319), .Z(n320) );
  GTECH_OR_NOT U222 ( .A(n330), .B(a[2]), .Z(n319) );
  GTECH_ADD_AB U223 ( .A(n329), .B(n330), .COUT(n317) );
  GTECH_NOT U224 ( .A(b[2]), .Z(n330) );
  GTECH_NOT U225 ( .A(a[2]), .Z(n329) );
  GTECH_AOI21 U226 ( .A(n326), .B(n334), .C(n328), .Z(n325) );
  GTECH_ADD_AB U227 ( .A(a[1]), .B(b[1]), .COUT(n328) );
  GTECH_NOT U228 ( .A(n383), .Z(n334) );
  GTECH_NOR2 U229 ( .A(a[0]), .B(b[0]), .Z(n383) );
  GTECH_OR2 U230 ( .A(b[1]), .B(a[1]), .Z(n326) );
  GTECH_OA21 U231 ( .A(a[7]), .B(n291), .C(n384), .Z(n380) );
  GTECH_AO21 U232 ( .A(n291), .B(a[7]), .C(b[7]), .Z(n384) );
  GTECH_OAI21 U233 ( .A(n301), .B(n293), .C(n295), .Z(n291) );
  GTECH_OR_NOT U234 ( .A(n385), .B(a[6]), .Z(n295) );
  GTECH_ADD_AB U235 ( .A(n300), .B(n385), .COUT(n293) );
  GTECH_NOT U236 ( .A(b[6]), .Z(n385) );
  GTECH_NOT U237 ( .A(a[6]), .Z(n300) );
  GTECH_AOI21 U238 ( .A(n386), .B(n303), .C(n305), .Z(n301) );
  GTECH_ADD_AB U239 ( .A(b[5]), .B(a[5]), .COUT(n305) );
  GTECH_OR2 U240 ( .A(b[5]), .B(a[5]), .Z(n303) );
  GTECH_OR2 U241 ( .A(b[4]), .B(a[4]), .Z(n386) );
  GTECH_XOR2 U242 ( .A(a[4]), .B(b[4]), .Z(n311) );
  GTECH_AOI21 U243 ( .A(n363), .B(a[11]), .C(n387), .Z(n379) );
  GTECH_OA21 U244 ( .A(a[11]), .B(n363), .C(b[11]), .Z(n387) );
  GTECH_OAI21 U245 ( .A(n372), .B(n365), .C(n367), .Z(n363) );
  GTECH_OR_NOT U246 ( .A(n388), .B(a[10]), .Z(n367) );
  GTECH_ADD_AB U247 ( .A(n389), .B(n388), .COUT(n365) );
  GTECH_NOT U248 ( .A(b[10]), .Z(n388) );
  GTECH_NOT U249 ( .A(a[10]), .Z(n389) );
  GTECH_AOI2N2 U250 ( .A(a[9]), .B(b[9]), .C(n283), .D(n285), .Z(n372) );
  GTECH_NOT U251 ( .A(n374), .Z(n285) );
  GTECH_OR2 U252 ( .A(b[9]), .B(a[9]), .Z(n374) );
  GTECH_NOT U253 ( .A(n286), .Z(n378) );
  GTECH_NOR2 U254 ( .A(n283), .B(n284), .Z(n286) );
  GTECH_ADD_AB U255 ( .A(b[8]), .B(a[8]), .COUT(n284) );
  GTECH_NOR2 U256 ( .A(a[8]), .B(b[8]), .Z(n283) );
  GTECH_OR_NOT U257 ( .A(n351), .B(n357), .Z(n359) );
  GTECH_ADD_AB U258 ( .A(a[12]), .B(b[12]), .COUT(n351) );
  GTECH_AOI21 U259 ( .A(n344), .B(a[15]), .C(n390), .Z(n377) );
  GTECH_NOT U260 ( .A(n391), .Z(n390) );
  GTECH_OAI21 U261 ( .A(a[15]), .B(n344), .C(b[15]), .Z(n391) );
  GTECH_OAI21 U262 ( .A(n340), .B(n350), .C(n342), .Z(n344) );
  GTECH_OR_NOT U263 ( .A(n349), .B(a[14]), .Z(n342) );
  GTECH_OAI21 U264 ( .A(n352), .B(n357), .C(n353), .Z(n350) );
  GTECH_OR_NOT U265 ( .A(b[13]), .B(n392), .Z(n353) );
  GTECH_NOT U266 ( .A(a[13]), .Z(n392) );
  GTECH_OR2 U267 ( .A(a[12]), .B(b[12]), .Z(n357) );
  GTECH_ADD_AB U268 ( .A(b[13]), .B(a[13]), .COUT(n352) );
  GTECH_ADD_AB U269 ( .A(n393), .B(n349), .COUT(n340) );
  GTECH_NOT U270 ( .A(b[14]), .Z(n349) );
  GTECH_NOT U271 ( .A(a[14]), .Z(n393) );
endmodule

