
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_NAND2 U83 ( .A(n93), .B(n94), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI22 U86 ( .A(n98), .B(n99), .C(n100), .D(n101), .Z(n89) );
  GTECH_AND2 U87 ( .A(n98), .B(n99), .Z(n100) );
  GTECH_NOT U88 ( .A(n102), .Z(n98) );
  GTECH_NAND2 U89 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U90 ( .A(n103), .Z(n84) );
  GTECH_NAND2 U91 ( .A(n104), .B(n105), .Z(n103) );
  GTECH_XOR2 U92 ( .A(n105), .B(n104), .Z(N153) );
  GTECH_NOT U93 ( .A(n106), .Z(n104) );
  GTECH_XOR3 U94 ( .A(n107), .B(n93), .C(n95), .Z(n106) );
  GTECH_XOR3 U95 ( .A(n108), .B(n109), .C(n102), .Z(n95) );
  GTECH_OAI22 U96 ( .A(n110), .B(n111), .C(n112), .D(n113), .Z(n102) );
  GTECH_AND2 U97 ( .A(n110), .B(n111), .Z(n112) );
  GTECH_NOT U98 ( .A(n114), .Z(n110) );
  GTECH_NOT U99 ( .A(n101), .Z(n109) );
  GTECH_NAND2 U100 ( .A(I_b[7]), .B(I_a[6]), .Z(n101) );
  GTECH_NOT U101 ( .A(n99), .Z(n108) );
  GTECH_NAND2 U102 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U103 ( .A(n115), .B(n116), .C(n117), .COUT(n93) );
  GTECH_NOT U104 ( .A(n118), .Z(n117) );
  GTECH_XOR2 U105 ( .A(n119), .B(n120), .Z(n116) );
  GTECH_AND2 U106 ( .A(I_a[7]), .B(I_b[5]), .Z(n120) );
  GTECH_NOT U107 ( .A(n94), .Z(n107) );
  GTECH_NAND2 U108 ( .A(I_a[7]), .B(n121), .Z(n94) );
  GTECH_NOT U109 ( .A(n122), .Z(n105) );
  GTECH_NAND2 U110 ( .A(n123), .B(n124), .Z(n122) );
  GTECH_NOT U111 ( .A(n125), .Z(n124) );
  GTECH_XOR2 U112 ( .A(n125), .B(n126), .Z(N152) );
  GTECH_NOT U113 ( .A(n123), .Z(n126) );
  GTECH_XOR4 U114 ( .A(n127), .B(n119), .C(n115), .D(n118), .Z(n123) );
  GTECH_XOR3 U115 ( .A(n128), .B(n129), .C(n114), .Z(n118) );
  GTECH_OAI22 U116 ( .A(n130), .B(n131), .C(n132), .D(n133), .Z(n114) );
  GTECH_AND2 U117 ( .A(n130), .B(n131), .Z(n132) );
  GTECH_NOT U118 ( .A(n134), .Z(n130) );
  GTECH_NOT U119 ( .A(n113), .Z(n129) );
  GTECH_NAND2 U120 ( .A(I_b[7]), .B(I_a[5]), .Z(n113) );
  GTECH_NOT U121 ( .A(n111), .Z(n128) );
  GTECH_NAND2 U122 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_ADD_ABC U123 ( .A(n135), .B(n136), .C(n137), .COUT(n115) );
  GTECH_NOT U124 ( .A(n138), .Z(n137) );
  GTECH_XOR3 U125 ( .A(n139), .B(n140), .C(n141), .Z(n136) );
  GTECH_NOT U126 ( .A(n142), .Z(n139) );
  GTECH_NOT U127 ( .A(n121), .Z(n119) );
  GTECH_OAI22 U128 ( .A(n141), .B(n142), .C(n143), .D(n144), .Z(n121) );
  GTECH_AND2 U129 ( .A(n141), .B(n142), .Z(n143) );
  GTECH_NOT U130 ( .A(n145), .Z(n141) );
  GTECH_AND2 U131 ( .A(I_a[7]), .B(I_b[5]), .Z(n127) );
  GTECH_ADD_ABC U132 ( .A(n146), .B(n147), .C(n148), .COUT(n125) );
  GTECH_NOT U133 ( .A(n149), .Z(n148) );
  GTECH_AOI2N2 U134 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n147) );
  GTECH_OA21 U135 ( .A(n154), .B(n155), .C(n156), .Z(n146) );
  GTECH_AO21 U136 ( .A(n154), .B(n155), .C(n157), .Z(n156) );
  GTECH_XOR3 U137 ( .A(n158), .B(n149), .C(n159), .Z(N151) );
  GTECH_OA21 U138 ( .A(n154), .B(n155), .C(n160), .Z(n159) );
  GTECH_AO21 U139 ( .A(n154), .B(n155), .C(n157), .Z(n160) );
  GTECH_XOR2 U140 ( .A(n161), .B(n135), .Z(n149) );
  GTECH_ADD_ABC U141 ( .A(n162), .B(n163), .C(n164), .COUT(n135) );
  GTECH_NOT U142 ( .A(n165), .Z(n164) );
  GTECH_XOR3 U143 ( .A(n166), .B(n167), .C(n168), .Z(n163) );
  GTECH_XOR4 U144 ( .A(n140), .B(n145), .C(n142), .D(n138), .Z(n161) );
  GTECH_XOR3 U145 ( .A(n169), .B(n170), .C(n134), .Z(n138) );
  GTECH_OAI22 U146 ( .A(n171), .B(n172), .C(n173), .D(n174), .Z(n134) );
  GTECH_AND2 U147 ( .A(n171), .B(n172), .Z(n173) );
  GTECH_NOT U148 ( .A(n175), .Z(n171) );
  GTECH_NOT U149 ( .A(n133), .Z(n170) );
  GTECH_NAND2 U150 ( .A(I_b[7]), .B(I_a[4]), .Z(n133) );
  GTECH_NOT U151 ( .A(n131), .Z(n169) );
  GTECH_NAND2 U152 ( .A(I_b[6]), .B(I_a[5]), .Z(n131) );
  GTECH_NAND2 U153 ( .A(I_a[7]), .B(I_b[4]), .Z(n142) );
  GTECH_OAI22 U154 ( .A(n168), .B(n176), .C(n177), .D(n178), .Z(n145) );
  GTECH_AND2 U155 ( .A(n168), .B(n176), .Z(n177) );
  GTECH_NOT U156 ( .A(n179), .Z(n168) );
  GTECH_NOT U157 ( .A(n144), .Z(n140) );
  GTECH_NAND2 U158 ( .A(I_a[6]), .B(I_b[5]), .Z(n144) );
  GTECH_AOI2N2 U159 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n158) );
  GTECH_NOT U160 ( .A(I_a[7]), .Z(n153) );
  GTECH_XOR3 U161 ( .A(n154), .B(n180), .C(n157), .Z(N150) );
  GTECH_XOR2 U162 ( .A(n162), .B(n181), .Z(n157) );
  GTECH_XOR4 U163 ( .A(n167), .B(n179), .C(n165), .D(n166), .Z(n181) );
  GTECH_NOT U164 ( .A(n176), .Z(n166) );
  GTECH_NAND2 U165 ( .A(I_a[6]), .B(I_b[4]), .Z(n176) );
  GTECH_XOR3 U166 ( .A(n182), .B(n183), .C(n175), .Z(n165) );
  GTECH_OAI22 U167 ( .A(n184), .B(n185), .C(n186), .D(n187), .Z(n175) );
  GTECH_AND2 U168 ( .A(n184), .B(n185), .Z(n186) );
  GTECH_NOT U169 ( .A(n188), .Z(n184) );
  GTECH_NOT U170 ( .A(n174), .Z(n183) );
  GTECH_NAND2 U171 ( .A(I_b[7]), .B(I_a[3]), .Z(n174) );
  GTECH_NOT U172 ( .A(n172), .Z(n182) );
  GTECH_NAND2 U173 ( .A(I_b[6]), .B(I_a[4]), .Z(n172) );
  GTECH_OAI22 U174 ( .A(n189), .B(n190), .C(n191), .D(n192), .Z(n179) );
  GTECH_AND2 U175 ( .A(n189), .B(n190), .Z(n191) );
  GTECH_NOT U176 ( .A(n178), .Z(n167) );
  GTECH_NAND2 U177 ( .A(I_a[5]), .B(I_b[5]), .Z(n178) );
  GTECH_ADD_ABC U178 ( .A(n193), .B(n194), .C(n195), .COUT(n162) );
  GTECH_NOT U179 ( .A(n196), .Z(n195) );
  GTECH_XOR3 U180 ( .A(n197), .B(n198), .C(n189), .Z(n194) );
  GTECH_NOT U181 ( .A(n199), .Z(n189) );
  GTECH_NOT U182 ( .A(n155), .Z(n180) );
  GTECH_XOR2 U183 ( .A(n150), .B(n200), .Z(n155) );
  GTECH_NOT U184 ( .A(n151), .Z(n200) );
  GTECH_OAI2N2 U185 ( .A(n201), .B(n202), .C(n203), .D(n204), .Z(n151) );
  GTECH_NAND2 U186 ( .A(n201), .B(n202), .Z(n204) );
  GTECH_XOR2 U187 ( .A(n205), .B(n152), .Z(n150) );
  GTECH_OA21 U188 ( .A(n206), .B(n207), .C(n208), .Z(n152) );
  GTECH_AO21 U189 ( .A(n206), .B(n207), .C(n209), .Z(n208) );
  GTECH_NOT U190 ( .A(n210), .Z(n206) );
  GTECH_NAND2 U191 ( .A(I_a[7]), .B(I_b[3]), .Z(n205) );
  GTECH_OA21 U192 ( .A(n211), .B(n212), .C(n213), .Z(n154) );
  GTECH_AO21 U193 ( .A(n211), .B(n212), .C(n214), .Z(n213) );
  GTECH_XOR3 U194 ( .A(n211), .B(n215), .C(n214), .Z(N149) );
  GTECH_XOR2 U195 ( .A(n193), .B(n216), .Z(n214) );
  GTECH_XOR4 U196 ( .A(n198), .B(n199), .C(n196), .D(n197), .Z(n216) );
  GTECH_NOT U197 ( .A(n190), .Z(n197) );
  GTECH_NAND2 U198 ( .A(I_a[5]), .B(I_b[4]), .Z(n190) );
  GTECH_XOR3 U199 ( .A(n217), .B(n218), .C(n188), .Z(n196) );
  GTECH_AO21 U200 ( .A(n219), .B(n220), .C(n221), .Z(n188) );
  GTECH_NOT U201 ( .A(n222), .Z(n221) );
  GTECH_NOT U202 ( .A(n187), .Z(n218) );
  GTECH_NAND2 U203 ( .A(I_b[7]), .B(I_a[2]), .Z(n187) );
  GTECH_NOT U204 ( .A(n185), .Z(n217) );
  GTECH_NAND2 U205 ( .A(I_b[6]), .B(I_a[3]), .Z(n185) );
  GTECH_OAI22 U206 ( .A(n223), .B(n224), .C(n225), .D(n226), .Z(n199) );
  GTECH_AND2 U207 ( .A(n223), .B(n224), .Z(n225) );
  GTECH_NOT U208 ( .A(n192), .Z(n198) );
  GTECH_NAND2 U209 ( .A(I_b[5]), .B(I_a[4]), .Z(n192) );
  GTECH_ADD_ABC U210 ( .A(n227), .B(n228), .C(n229), .COUT(n193) );
  GTECH_XOR3 U211 ( .A(n230), .B(n231), .C(n223), .Z(n228) );
  GTECH_NOT U212 ( .A(n232), .Z(n223) );
  GTECH_NOT U213 ( .A(n224), .Z(n230) );
  GTECH_OA21 U214 ( .A(n233), .B(n234), .C(n235), .Z(n227) );
  GTECH_AO21 U215 ( .A(n233), .B(n234), .C(n236), .Z(n235) );
  GTECH_NOT U216 ( .A(n212), .Z(n215) );
  GTECH_XOR3 U217 ( .A(n237), .B(n201), .C(n203), .Z(n212) );
  GTECH_XOR3 U218 ( .A(n238), .B(n239), .C(n210), .Z(n203) );
  GTECH_OAI22 U219 ( .A(n240), .B(n241), .C(n242), .D(n243), .Z(n210) );
  GTECH_AND2 U220 ( .A(n240), .B(n241), .Z(n242) );
  GTECH_NOT U221 ( .A(n244), .Z(n240) );
  GTECH_NOT U222 ( .A(n209), .Z(n239) );
  GTECH_NAND2 U223 ( .A(I_a[6]), .B(I_b[3]), .Z(n209) );
  GTECH_NOT U224 ( .A(n207), .Z(n238) );
  GTECH_NAND2 U225 ( .A(I_a[7]), .B(I_b[2]), .Z(n207) );
  GTECH_ADD_ABC U226 ( .A(n245), .B(n246), .C(n247), .COUT(n201) );
  GTECH_XOR2 U227 ( .A(n248), .B(n249), .Z(n246) );
  GTECH_AND2 U228 ( .A(I_a[7]), .B(I_b[1]), .Z(n249) );
  GTECH_NOT U229 ( .A(n202), .Z(n237) );
  GTECH_NAND2 U230 ( .A(I_a[7]), .B(n250), .Z(n202) );
  GTECH_ADD_ABC U231 ( .A(n251), .B(n252), .C(n253), .COUT(n211) );
  GTECH_XOR3 U232 ( .A(n245), .B(n254), .C(n247), .Z(n252) );
  GTECH_NOT U233 ( .A(n255), .Z(n247) );
  GTECH_XOR2 U234 ( .A(n251), .B(n256), .Z(N148) );
  GTECH_XOR4 U235 ( .A(n254), .B(n255), .C(n253), .D(n245), .Z(n256) );
  GTECH_ADD_ABC U236 ( .A(n257), .B(n258), .C(n259), .COUT(n245) );
  GTECH_XOR3 U237 ( .A(n260), .B(n261), .C(n262), .Z(n258) );
  GTECH_XOR2 U238 ( .A(n263), .B(n264), .Z(n253) );
  GTECH_OA21 U239 ( .A(n233), .B(n234), .C(n265), .Z(n264) );
  GTECH_AO21 U240 ( .A(n233), .B(n234), .C(n236), .Z(n265) );
  GTECH_XOR4 U241 ( .A(n231), .B(n232), .C(n224), .D(n229), .Z(n263) );
  GTECH_XOR3 U242 ( .A(n220), .B(n219), .C(n222), .Z(n229) );
  GTECH_NAND3 U243 ( .A(I_b[6]), .B(I_a[1]), .C(n266), .Z(n222) );
  GTECH_NOT U244 ( .A(n267), .Z(n219) );
  GTECH_NAND2 U245 ( .A(I_b[7]), .B(I_a[1]), .Z(n267) );
  GTECH_NOT U246 ( .A(n268), .Z(n220) );
  GTECH_NAND2 U247 ( .A(I_b[6]), .B(I_a[2]), .Z(n268) );
  GTECH_NAND2 U248 ( .A(I_b[4]), .B(I_a[4]), .Z(n224) );
  GTECH_OAI22 U249 ( .A(n269), .B(n270), .C(n271), .D(n272), .Z(n232) );
  GTECH_AND2 U250 ( .A(n269), .B(n270), .Z(n271) );
  GTECH_NOT U251 ( .A(n273), .Z(n269) );
  GTECH_NOT U252 ( .A(n226), .Z(n231) );
  GTECH_NAND2 U253 ( .A(I_b[5]), .B(I_a[3]), .Z(n226) );
  GTECH_XOR3 U254 ( .A(n274), .B(n275), .C(n244), .Z(n255) );
  GTECH_OAI22 U255 ( .A(n276), .B(n277), .C(n278), .D(n279), .Z(n244) );
  GTECH_AND2 U256 ( .A(n276), .B(n277), .Z(n278) );
  GTECH_NOT U257 ( .A(n280), .Z(n276) );
  GTECH_NOT U258 ( .A(n243), .Z(n275) );
  GTECH_NAND2 U259 ( .A(I_a[5]), .B(I_b[3]), .Z(n243) );
  GTECH_NOT U260 ( .A(n241), .Z(n274) );
  GTECH_NAND2 U261 ( .A(I_a[6]), .B(I_b[2]), .Z(n241) );
  GTECH_XOR2 U262 ( .A(n281), .B(n248), .Z(n254) );
  GTECH_NOT U263 ( .A(n250), .Z(n248) );
  GTECH_OAI22 U264 ( .A(n262), .B(n282), .C(n283), .D(n284), .Z(n250) );
  GTECH_AND2 U265 ( .A(n262), .B(n282), .Z(n283) );
  GTECH_NOT U266 ( .A(n285), .Z(n262) );
  GTECH_AND2 U267 ( .A(I_a[7]), .B(I_b[1]), .Z(n281) );
  GTECH_ADD_ABC U268 ( .A(n286), .B(n287), .C(n288), .COUT(n251) );
  GTECH_NOT U269 ( .A(n289), .Z(n288) );
  GTECH_XOR3 U270 ( .A(n257), .B(n290), .C(n259), .Z(n287) );
  GTECH_NOT U271 ( .A(n291), .Z(n259) );
  GTECH_NOT U272 ( .A(n292), .Z(n290) );
  GTECH_XOR2 U273 ( .A(n293), .B(n286), .Z(N147) );
  GTECH_ADD_ABC U274 ( .A(n294), .B(n295), .C(n296), .COUT(n286) );
  GTECH_XOR3 U275 ( .A(n297), .B(n298), .C(n299), .Z(n295) );
  GTECH_OA21 U276 ( .A(n300), .B(n301), .C(n302), .Z(n294) );
  GTECH_AO21 U277 ( .A(n300), .B(n301), .C(n303), .Z(n302) );
  GTECH_XOR4 U278 ( .A(n291), .B(n257), .C(n292), .D(n289), .Z(n293) );
  GTECH_XOR3 U279 ( .A(n304), .B(n234), .C(n233), .Z(n289) );
  GTECH_XOR2 U280 ( .A(n305), .B(n266), .Z(n233) );
  GTECH_NOT U281 ( .A(n306), .Z(n266) );
  GTECH_NAND2 U282 ( .A(I_b[7]), .B(I_a[0]), .Z(n306) );
  GTECH_NAND2 U283 ( .A(I_b[6]), .B(I_a[1]), .Z(n305) );
  GTECH_NOT U284 ( .A(n307), .Z(n234) );
  GTECH_XOR3 U285 ( .A(n308), .B(n309), .C(n273), .Z(n307) );
  GTECH_AO21 U286 ( .A(n310), .B(n311), .C(n312), .Z(n273) );
  GTECH_NOT U287 ( .A(n313), .Z(n312) );
  GTECH_NOT U288 ( .A(n272), .Z(n309) );
  GTECH_NAND2 U289 ( .A(I_b[5]), .B(I_a[2]), .Z(n272) );
  GTECH_NOT U290 ( .A(n270), .Z(n308) );
  GTECH_NAND2 U291 ( .A(I_b[4]), .B(I_a[3]), .Z(n270) );
  GTECH_NOT U292 ( .A(n236), .Z(n304) );
  GTECH_NAND3 U293 ( .A(I_a[0]), .B(n314), .C(I_b[6]), .Z(n236) );
  GTECH_NOT U294 ( .A(n315), .Z(n314) );
  GTECH_XOR3 U295 ( .A(n260), .B(n261), .C(n285), .Z(n292) );
  GTECH_OAI22 U296 ( .A(n316), .B(n317), .C(n318), .D(n319), .Z(n285) );
  GTECH_AND2 U297 ( .A(n316), .B(n317), .Z(n318) );
  GTECH_NOT U298 ( .A(n284), .Z(n261) );
  GTECH_NAND2 U299 ( .A(I_a[6]), .B(I_b[1]), .Z(n284) );
  GTECH_NOT U300 ( .A(n282), .Z(n260) );
  GTECH_NAND2 U301 ( .A(I_a[7]), .B(I_b[0]), .Z(n282) );
  GTECH_ADD_ABC U302 ( .A(n297), .B(n320), .C(n299), .COUT(n257) );
  GTECH_NOT U303 ( .A(n321), .Z(n299) );
  GTECH_XOR3 U304 ( .A(n322), .B(n323), .C(n316), .Z(n320) );
  GTECH_NOT U305 ( .A(n324), .Z(n316) );
  GTECH_XOR3 U306 ( .A(n325), .B(n326), .C(n280), .Z(n291) );
  GTECH_OAI22 U307 ( .A(n327), .B(n328), .C(n329), .D(n330), .Z(n280) );
  GTECH_AND2 U308 ( .A(n327), .B(n328), .Z(n329) );
  GTECH_NOT U309 ( .A(n331), .Z(n327) );
  GTECH_NOT U310 ( .A(n279), .Z(n326) );
  GTECH_NAND2 U311 ( .A(I_b[3]), .B(I_a[4]), .Z(n279) );
  GTECH_NOT U312 ( .A(n277), .Z(n325) );
  GTECH_NAND2 U313 ( .A(I_a[5]), .B(I_b[2]), .Z(n277) );
  GTECH_XOR2 U314 ( .A(n332), .B(n333), .Z(N146) );
  GTECH_XOR4 U315 ( .A(n298), .B(n321), .C(n296), .D(n297), .Z(n333) );
  GTECH_ADD_ABC U316 ( .A(n334), .B(n335), .C(n336), .COUT(n297) );
  GTECH_NOT U317 ( .A(n337), .Z(n336) );
  GTECH_XOR3 U318 ( .A(n338), .B(n339), .C(n340), .Z(n335) );
  GTECH_XOR2 U319 ( .A(n315), .B(n341), .Z(n296) );
  GTECH_AND2 U320 ( .A(I_b[6]), .B(I_a[0]), .Z(n341) );
  GTECH_XOR3 U321 ( .A(n311), .B(n310), .C(n313), .Z(n315) );
  GTECH_NAND3 U322 ( .A(I_b[4]), .B(I_a[1]), .C(n342), .Z(n313) );
  GTECH_NOT U323 ( .A(n343), .Z(n310) );
  GTECH_NAND2 U324 ( .A(I_b[5]), .B(I_a[1]), .Z(n343) );
  GTECH_NOT U325 ( .A(n344), .Z(n311) );
  GTECH_NAND2 U326 ( .A(I_b[4]), .B(I_a[2]), .Z(n344) );
  GTECH_XOR3 U327 ( .A(n345), .B(n346), .C(n331), .Z(n321) );
  GTECH_OAI22 U328 ( .A(n347), .B(n348), .C(n349), .D(n350), .Z(n331) );
  GTECH_AND2 U329 ( .A(n347), .B(n348), .Z(n349) );
  GTECH_NOT U330 ( .A(n351), .Z(n347) );
  GTECH_NOT U331 ( .A(n330), .Z(n346) );
  GTECH_NAND2 U332 ( .A(I_b[3]), .B(I_a[3]), .Z(n330) );
  GTECH_NOT U333 ( .A(n328), .Z(n345) );
  GTECH_NAND2 U334 ( .A(I_b[2]), .B(I_a[4]), .Z(n328) );
  GTECH_NOT U335 ( .A(n352), .Z(n298) );
  GTECH_XOR3 U336 ( .A(n322), .B(n323), .C(n324), .Z(n352) );
  GTECH_OAI22 U337 ( .A(n340), .B(n353), .C(n354), .D(n355), .Z(n324) );
  GTECH_AND2 U338 ( .A(n340), .B(n353), .Z(n354) );
  GTECH_NOT U339 ( .A(n356), .Z(n340) );
  GTECH_NOT U340 ( .A(n319), .Z(n323) );
  GTECH_NAND2 U341 ( .A(I_a[5]), .B(I_b[1]), .Z(n319) );
  GTECH_NOT U342 ( .A(n317), .Z(n322) );
  GTECH_NAND2 U343 ( .A(I_a[6]), .B(I_b[0]), .Z(n317) );
  GTECH_OA21 U344 ( .A(n300), .B(n301), .C(n357), .Z(n332) );
  GTECH_AO21 U345 ( .A(n300), .B(n301), .C(n303), .Z(n357) );
  GTECH_XOR3 U346 ( .A(n358), .B(n301), .C(n300), .Z(N145) );
  GTECH_XOR2 U347 ( .A(n359), .B(n342), .Z(n300) );
  GTECH_NOT U348 ( .A(n360), .Z(n342) );
  GTECH_NAND2 U349 ( .A(I_b[5]), .B(I_a[0]), .Z(n360) );
  GTECH_NAND2 U350 ( .A(I_b[4]), .B(I_a[1]), .Z(n359) );
  GTECH_XOR2 U351 ( .A(n334), .B(n361), .Z(n301) );
  GTECH_XOR4 U352 ( .A(n339), .B(n356), .C(n337), .D(n338), .Z(n361) );
  GTECH_NOT U353 ( .A(n353), .Z(n338) );
  GTECH_NAND2 U354 ( .A(I_a[5]), .B(I_b[0]), .Z(n353) );
  GTECH_XOR3 U355 ( .A(n362), .B(n363), .C(n351), .Z(n337) );
  GTECH_AO21 U356 ( .A(n364), .B(n365), .C(n366), .Z(n351) );
  GTECH_NOT U357 ( .A(n367), .Z(n366) );
  GTECH_NOT U358 ( .A(n350), .Z(n363) );
  GTECH_NAND2 U359 ( .A(I_b[3]), .B(I_a[2]), .Z(n350) );
  GTECH_NOT U360 ( .A(n348), .Z(n362) );
  GTECH_NAND2 U361 ( .A(I_b[2]), .B(I_a[3]), .Z(n348) );
  GTECH_OAI22 U362 ( .A(n368), .B(n369), .C(n370), .D(n371), .Z(n356) );
  GTECH_AND2 U363 ( .A(n368), .B(n369), .Z(n370) );
  GTECH_NOT U364 ( .A(n355), .Z(n339) );
  GTECH_NAND2 U365 ( .A(I_a[4]), .B(I_b[1]), .Z(n355) );
  GTECH_ADD_ABC U366 ( .A(n372), .B(n373), .C(n374), .COUT(n334) );
  GTECH_XOR3 U367 ( .A(n375), .B(n376), .C(n368), .Z(n373) );
  GTECH_NOT U368 ( .A(n377), .Z(n368) );
  GTECH_OA21 U369 ( .A(n378), .B(n379), .C(n380), .Z(n372) );
  GTECH_AO21 U370 ( .A(n378), .B(n379), .C(n381), .Z(n380) );
  GTECH_NOT U371 ( .A(n303), .Z(n358) );
  GTECH_NAND3 U372 ( .A(I_a[0]), .B(n382), .C(I_b[4]), .Z(n303) );
  GTECH_XOR2 U373 ( .A(n383), .B(n382), .Z(N144) );
  GTECH_XOR2 U374 ( .A(n384), .B(n385), .Z(n382) );
  GTECH_XOR4 U375 ( .A(n376), .B(n377), .C(n374), .D(n375), .Z(n385) );
  GTECH_NOT U376 ( .A(n369), .Z(n375) );
  GTECH_NAND2 U377 ( .A(I_a[4]), .B(I_b[0]), .Z(n369) );
  GTECH_XOR3 U378 ( .A(n365), .B(n364), .C(n367), .Z(n374) );
  GTECH_NAND3 U379 ( .A(I_b[2]), .B(I_a[1]), .C(n386), .Z(n367) );
  GTECH_NOT U380 ( .A(n387), .Z(n364) );
  GTECH_NAND2 U381 ( .A(I_b[3]), .B(I_a[1]), .Z(n387) );
  GTECH_NOT U382 ( .A(n388), .Z(n365) );
  GTECH_NAND2 U383 ( .A(I_b[2]), .B(I_a[2]), .Z(n388) );
  GTECH_OAI22 U384 ( .A(n389), .B(n390), .C(n391), .D(n392), .Z(n377) );
  GTECH_AND2 U385 ( .A(n389), .B(n390), .Z(n391) );
  GTECH_NOT U386 ( .A(n393), .Z(n389) );
  GTECH_NOT U387 ( .A(n371), .Z(n376) );
  GTECH_NAND2 U388 ( .A(I_a[3]), .B(I_b[1]), .Z(n371) );
  GTECH_OA21 U389 ( .A(n378), .B(n379), .C(n394), .Z(n384) );
  GTECH_AO21 U390 ( .A(n378), .B(n379), .C(n381), .Z(n394) );
  GTECH_AND2 U391 ( .A(I_b[4]), .B(I_a[0]), .Z(n383) );
  GTECH_XOR3 U392 ( .A(n395), .B(n379), .C(n378), .Z(N143) );
  GTECH_XOR2 U393 ( .A(n396), .B(n386), .Z(n378) );
  GTECH_NOT U394 ( .A(n397), .Z(n386) );
  GTECH_NAND2 U395 ( .A(I_b[3]), .B(I_a[0]), .Z(n397) );
  GTECH_NAND2 U396 ( .A(I_b[2]), .B(I_a[1]), .Z(n396) );
  GTECH_NOT U397 ( .A(n398), .Z(n379) );
  GTECH_XOR3 U398 ( .A(n399), .B(n400), .C(n393), .Z(n398) );
  GTECH_AO21 U399 ( .A(n401), .B(n402), .C(n403), .Z(n393) );
  GTECH_NOT U400 ( .A(n404), .Z(n403) );
  GTECH_NOT U401 ( .A(n392), .Z(n400) );
  GTECH_NAND2 U402 ( .A(I_b[1]), .B(I_a[2]), .Z(n392) );
  GTECH_NOT U403 ( .A(n390), .Z(n399) );
  GTECH_NAND2 U404 ( .A(I_b[0]), .B(I_a[3]), .Z(n390) );
  GTECH_NOT U405 ( .A(n381), .Z(n395) );
  GTECH_NAND3 U406 ( .A(I_a[0]), .B(n405), .C(I_b[2]), .Z(n381) );
  GTECH_XOR2 U407 ( .A(n406), .B(n405), .Z(N142) );
  GTECH_NOT U408 ( .A(n407), .Z(n405) );
  GTECH_XOR3 U409 ( .A(n401), .B(n402), .C(n404), .Z(n407) );
  GTECH_NAND3 U410 ( .A(n408), .B(I_b[0]), .C(I_a[1]), .Z(n404) );
  GTECH_NOT U411 ( .A(n409), .Z(n402) );
  GTECH_NAND2 U412 ( .A(I_a[1]), .B(I_b[1]), .Z(n409) );
  GTECH_NOT U413 ( .A(n410), .Z(n401) );
  GTECH_NAND2 U414 ( .A(I_b[0]), .B(I_a[2]), .Z(n410) );
  GTECH_AND2 U415 ( .A(I_b[2]), .B(I_a[0]), .Z(n406) );
  GTECH_XOR2 U416 ( .A(n408), .B(n411), .Z(N141) );
  GTECH_AND2 U417 ( .A(I_a[1]), .B(I_b[0]), .Z(n411) );
  GTECH_NOT U418 ( .A(n412), .Z(n408) );
  GTECH_NAND2 U419 ( .A(I_a[0]), .B(I_b[1]), .Z(n412) );
  GTECH_AND2 U420 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

