
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374;

  GTECH_MUX2 U131 ( .A(n270), .B(n271), .S(n272), .Z(sum[9]) );
  GTECH_OA21 U132 ( .A(n273), .B(n274), .C(n275), .Z(n272) );
  GTECH_OAI21 U133 ( .A(a[8]), .B(n276), .C(b[8]), .Z(n275) );
  GTECH_NOT U134 ( .A(a[8]), .Z(n274) );
  GTECH_XOR2 U135 ( .A(b[9]), .B(a[9]), .Z(n271) );
  GTECH_OR_NOT U136 ( .A(n277), .B(n278), .Z(n270) );
  GTECH_OAI21 U137 ( .A(n273), .B(n279), .C(n280), .Z(sum[8]) );
  GTECH_MUX2 U138 ( .A(n281), .B(n282), .S(n283), .Z(sum[7]) );
  GTECH_XOR2 U139 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_XOR2 U140 ( .A(n286), .B(n285), .Z(n281) );
  GTECH_XOR2 U141 ( .A(a[7]), .B(b[7]), .Z(n285) );
  GTECH_OA21 U142 ( .A(n287), .B(n288), .C(n289), .Z(n286) );
  GTECH_MUX2 U143 ( .A(n290), .B(n291), .S(n283), .Z(sum[6]) );
  GTECH_XNOR2 U144 ( .A(n292), .B(n293), .Z(n291) );
  GTECH_XNOR2 U145 ( .A(n292), .B(n288), .Z(n290) );
  GTECH_OAI21 U146 ( .A(n294), .B(n295), .C(n296), .Z(n288) );
  GTECH_OAI21 U147 ( .A(a[6]), .B(b[6]), .C(n297), .Z(n292) );
  GTECH_NOT U148 ( .A(n287), .Z(n297) );
  GTECH_MUX2 U149 ( .A(n298), .B(n299), .S(n300), .Z(sum[5]) );
  GTECH_AND_NOT U150 ( .A(n296), .B(n294), .Z(n300) );
  GTECH_OAI2N2 U151 ( .A(b[4]), .B(a[4]), .C(n295), .D(n301), .Z(n299) );
  GTECH_NOT U152 ( .A(n283), .Z(n301) );
  GTECH_NAND2 U153 ( .A(b[4]), .B(a[4]), .Z(n295) );
  GTECH_ADD_ABC U154 ( .A(n283), .B(a[4]), .C(b[4]), .COUT(n298) );
  GTECH_XOR2 U155 ( .A(n283), .B(n302), .Z(sum[4]) );
  GTECH_MUX2 U156 ( .A(n303), .B(n304), .S(cin), .Z(sum[3]) );
  GTECH_XOR2 U157 ( .A(n305), .B(n306), .Z(n304) );
  GTECH_XOR2 U158 ( .A(n307), .B(n306), .Z(n303) );
  GTECH_XOR2 U159 ( .A(a[3]), .B(b[3]), .Z(n306) );
  GTECH_OA21 U160 ( .A(n308), .B(n309), .C(n310), .Z(n307) );
  GTECH_MUX2 U161 ( .A(n311), .B(n312), .S(cin), .Z(sum[2]) );
  GTECH_XOR2 U162 ( .A(n313), .B(n314), .Z(n312) );
  GTECH_XOR2 U163 ( .A(n309), .B(n313), .Z(n311) );
  GTECH_OA21 U164 ( .A(a[2]), .B(b[2]), .C(n315), .Z(n313) );
  GTECH_NOT U165 ( .A(n308), .Z(n315) );
  GTECH_OAI21 U166 ( .A(n316), .B(n317), .C(n318), .Z(n309) );
  GTECH_MUX2 U167 ( .A(n319), .B(n320), .S(n321), .Z(sum[1]) );
  GTECH_AND_NOT U168 ( .A(n318), .B(n316), .Z(n321) );
  GTECH_OAI21 U169 ( .A(cin), .B(n322), .C(n323), .Z(n320) );
  GTECH_NOT U170 ( .A(n317), .Z(n322) );
  GTECH_OAI21 U171 ( .A(n324), .B(n325), .C(n317), .Z(n319) );
  GTECH_MUX2 U172 ( .A(n326), .B(n327), .S(n328), .Z(sum[15]) );
  GTECH_XNOR2 U173 ( .A(n329), .B(n330), .Z(n327) );
  GTECH_XNOR2 U174 ( .A(n331), .B(n330), .Z(n326) );
  GTECH_XNOR2 U175 ( .A(a[15]), .B(b[15]), .Z(n330) );
  GTECH_OA21 U176 ( .A(n332), .B(n333), .C(n334), .Z(n331) );
  GTECH_MUX2 U177 ( .A(n335), .B(n336), .S(n328), .Z(sum[14]) );
  GTECH_XOR2 U178 ( .A(n337), .B(n338), .Z(n336) );
  GTECH_XOR2 U179 ( .A(n337), .B(n333), .Z(n335) );
  GTECH_OA21 U180 ( .A(n339), .B(n340), .C(n341), .Z(n333) );
  GTECH_OA21 U181 ( .A(a[14]), .B(b[14]), .C(n342), .Z(n337) );
  GTECH_NOT U182 ( .A(n332), .Z(n342) );
  GTECH_MUX2 U183 ( .A(n343), .B(n344), .S(n328), .Z(sum[13]) );
  GTECH_XOR2 U184 ( .A(n345), .B(n346), .Z(n344) );
  GTECH_XOR2 U185 ( .A(n345), .B(n340), .Z(n343) );
  GTECH_OA21 U186 ( .A(a[13]), .B(b[13]), .C(n347), .Z(n345) );
  GTECH_NOT U187 ( .A(n339), .Z(n347) );
  GTECH_NAND2 U188 ( .A(n348), .B(n349), .Z(sum[12]) );
  GTECH_OAI21 U189 ( .A(n340), .B(n350), .C(n328), .Z(n348) );
  GTECH_MUX2 U190 ( .A(n351), .B(n352), .S(n273), .Z(sum[11]) );
  GTECH_XOR2 U191 ( .A(n353), .B(n354), .Z(n352) );
  GTECH_OA21 U192 ( .A(n355), .B(n356), .C(n357), .Z(n353) );
  GTECH_XOR2 U193 ( .A(n358), .B(n354), .Z(n351) );
  GTECH_XOR2 U194 ( .A(a[11]), .B(b[11]), .Z(n354) );
  GTECH_MUX2 U195 ( .A(n359), .B(n360), .S(n273), .Z(sum[10]) );
  GTECH_XNOR2 U196 ( .A(n361), .B(n356), .Z(n360) );
  GTECH_OR_NOT U197 ( .A(n277), .B(n362), .Z(n356) );
  GTECH_NAND3 U198 ( .A(b[8]), .B(n278), .C(a[8]), .Z(n362) );
  GTECH_XNOR2 U199 ( .A(n361), .B(n363), .Z(n359) );
  GTECH_OAI21 U200 ( .A(a[10]), .B(b[10]), .C(n364), .Z(n361) );
  GTECH_NOT U201 ( .A(n355), .Z(n364) );
  GTECH_XNOR2 U202 ( .A(n325), .B(n365), .Z(sum[0]) );
  GTECH_NOT U203 ( .A(cin), .Z(n325) );
  GTECH_NAND2 U204 ( .A(n366), .B(n349), .Z(cout) );
  GTECH_OR3 U205 ( .A(n340), .B(n350), .C(n328), .Z(n349) );
  GTECH_AND2 U206 ( .A(b[12]), .B(a[12]), .Z(n340) );
  GTECH_NAND2 U207 ( .A(n367), .B(n328), .Z(n366) );
  GTECH_NAND2 U208 ( .A(n368), .B(n280), .Z(n328) );
  GTECH_OR_NOT U209 ( .A(n276), .B(n279), .Z(n280) );
  GTECH_XOR2 U210 ( .A(a[8]), .B(b[8]), .Z(n279) );
  GTECH_OR_NOT U211 ( .A(n273), .B(n369), .Z(n368) );
  GTECH_ADD_ABC U212 ( .A(a[11]), .B(n358), .C(b[11]), .COUT(n369) );
  GTECH_OA21 U213 ( .A(n355), .B(n363), .C(n357), .Z(n358) );
  GTECH_OR2 U214 ( .A(b[10]), .B(a[10]), .Z(n357) );
  GTECH_OR_NOT U215 ( .A(n277), .B(n370), .Z(n363) );
  GTECH_OAI21 U216 ( .A(b[8]), .B(a[8]), .C(n278), .Z(n370) );
  GTECH_OR2 U217 ( .A(a[9]), .B(b[9]), .Z(n278) );
  GTECH_AND2 U218 ( .A(b[9]), .B(a[9]), .Z(n277) );
  GTECH_AND2 U219 ( .A(b[10]), .B(a[10]), .Z(n355) );
  GTECH_NOT U220 ( .A(n276), .Z(n273) );
  GTECH_MUX2 U221 ( .A(n302), .B(n371), .S(n283), .Z(n276) );
  GTECH_MUX2 U222 ( .A(n365), .B(n372), .S(cin), .Z(n283) );
  GTECH_ADD_ABC U223 ( .A(n305), .B(a[3]), .C(b[3]), .COUT(n372) );
  GTECH_OA21 U224 ( .A(n308), .B(n314), .C(n310), .Z(n305) );
  GTECH_OR2 U225 ( .A(b[2]), .B(a[2]), .Z(n310) );
  GTECH_OAI21 U226 ( .A(n324), .B(n316), .C(n318), .Z(n314) );
  GTECH_NAND2 U227 ( .A(b[1]), .B(a[1]), .Z(n318) );
  GTECH_NOR2 U228 ( .A(a[1]), .B(b[1]), .Z(n316) );
  GTECH_AND2 U229 ( .A(b[2]), .B(a[2]), .Z(n308) );
  GTECH_AND2 U230 ( .A(n323), .B(n317), .Z(n365) );
  GTECH_NAND2 U231 ( .A(b[0]), .B(a[0]), .Z(n317) );
  GTECH_NOT U232 ( .A(n324), .Z(n323) );
  GTECH_NOR2 U233 ( .A(b[0]), .B(a[0]), .Z(n324) );
  GTECH_ADD_ABC U234 ( .A(a[7]), .B(n284), .C(b[7]), .COUT(n371) );
  GTECH_OA21 U235 ( .A(n287), .B(n293), .C(n289), .Z(n284) );
  GTECH_OR2 U236 ( .A(b[6]), .B(a[6]), .Z(n289) );
  GTECH_NAND2 U237 ( .A(n373), .B(n296), .Z(n293) );
  GTECH_NAND2 U238 ( .A(b[5]), .B(a[5]), .Z(n296) );
  GTECH_OAI21 U239 ( .A(b[4]), .B(a[4]), .C(n374), .Z(n373) );
  GTECH_NOT U240 ( .A(n294), .Z(n374) );
  GTECH_NOR2 U241 ( .A(a[5]), .B(b[5]), .Z(n294) );
  GTECH_AND2 U242 ( .A(b[6]), .B(a[6]), .Z(n287) );
  GTECH_XOR2 U243 ( .A(a[4]), .B(b[4]), .Z(n302) );
  GTECH_ADD_ABC U244 ( .A(a[15]), .B(n329), .C(b[15]), .COUT(n367) );
  GTECH_OA21 U245 ( .A(n332), .B(n338), .C(n334), .Z(n329) );
  GTECH_OR2 U246 ( .A(b[14]), .B(a[14]), .Z(n334) );
  GTECH_OA21 U247 ( .A(n339), .B(n346), .C(n341), .Z(n338) );
  GTECH_OR2 U248 ( .A(b[13]), .B(a[13]), .Z(n341) );
  GTECH_NOT U249 ( .A(n350), .Z(n346) );
  GTECH_NOR2 U250 ( .A(a[12]), .B(b[12]), .Z(n350) );
  GTECH_AND2 U251 ( .A(b[13]), .B(a[13]), .Z(n339) );
  GTECH_AND2 U252 ( .A(b[14]), .B(a[14]), .Z(n332) );
endmodule

