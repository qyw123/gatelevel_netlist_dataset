
module clock_12h ( clk, reset, ena, pm, hh, mm, ss );
  output [7:0] hh;
  output [7:0] mm;
  output [7:0] ss;
  input clk, reset, ena;
  output pm;
  wire   N22, N23, N24, N25, N26, N39, N40, N41, N42, N43, N55, N56, N57, N58,
         N59, N71, N72, N73, N74, N75, N88, N89, N90, N91, N92, N110, N112,
         N114, N115, N116, N121, N122, n3, n4, n5, n6, n7, n8, n9, n84, n109,
         n110, n111, n112, n113, n114, n115, n116, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217;

  GTECH_FJK1S ss_ones_reg_0_ ( .J(n84), .K(n84), .TI(N22), .TE(N25), .CP(clk), 
        .Q(ss[0]) );
  GTECH_FJK1S ss_ones_reg_2_ ( .J(n84), .K(n84), .TI(N24), .TE(N25), .CP(clk), 
        .Q(ss[2]) );
  GTECH_FJK1S ss_ones_reg_3_ ( .J(n84), .K(n84), .TI(N26), .TE(N25), .CP(clk), 
        .Q(ss[3]) );
  GTECH_FJK1S ss_ones_reg_1_ ( .J(n84), .K(n84), .TI(N23), .TE(N25), .CP(clk), 
        .Q(ss[1]) );
  GTECH_FJK1S ss_tens_reg_0_ ( .J(n84), .K(n84), .TI(N39), .TE(N42), .CP(clk), 
        .Q(ss[4]) );
  GTECH_FJK1S ss_tens_reg_2_ ( .J(n84), .K(n84), .TI(N41), .TE(N42), .CP(clk), 
        .Q(ss[6]) );
  GTECH_FJK1S ss_tens_reg_3_ ( .J(n84), .K(n84), .TI(N43), .TE(N42), .CP(clk), 
        .Q(ss[7]) );
  GTECH_FJK1S ss_tens_reg_1_ ( .J(n84), .K(n84), .TI(N40), .TE(N42), .CP(clk), 
        .Q(ss[5]) );
  GTECH_FJK1S mm_ones_reg_0_ ( .J(n84), .K(n84), .TI(N55), .TE(N58), .CP(clk), 
        .Q(mm[0]), .QN(n114) );
  GTECH_FJK1S mm_ones_reg_2_ ( .J(n84), .K(n84), .TI(N57), .TE(N58), .CP(clk), 
        .Q(mm[2]), .QN(n116) );
  GTECH_FJK1S mm_ones_reg_3_ ( .J(n84), .K(n84), .TI(N59), .TE(N58), .CP(clk), 
        .Q(mm[3]), .QN(n113) );
  GTECH_FJK1S mm_ones_reg_1_ ( .J(n84), .K(n84), .TI(N56), .TE(N58), .CP(clk), 
        .Q(mm[1]), .QN(n115) );
  GTECH_FJK1S mm_tens_reg_0_ ( .J(n84), .K(n84), .TI(N71), .TE(N74), .CP(clk), 
        .Q(mm[4]), .QN(n3) );
  GTECH_FJK1S mm_tens_reg_2_ ( .J(n84), .K(n84), .TI(N73), .TE(N74), .CP(clk), 
        .Q(mm[6]), .QN(n111) );
  GTECH_FJK1S mm_tens_reg_3_ ( .J(n84), .K(n84), .TI(N75), .TE(N74), .CP(clk), 
        .Q(mm[7]), .QN(n110) );
  GTECH_FJK1S mm_tens_reg_1_ ( .J(n84), .K(n84), .TI(N72), .TE(N74), .CP(clk), 
        .Q(mm[5]), .QN(n112) );
  GTECH_FJK1S hh_tens_reg_0_ ( .J(n84), .K(n84), .TI(N110), .TE(N115), .CP(clk), .Q(hh[4]), .QN(n4) );
  GTECH_FJK1S hh_tens_reg_2_ ( .J(n84), .K(n84), .TI(N114), .TE(N115), .CP(clk), .Q(hh[6]), .QN(n5) );
  GTECH_FJK1S hh_tens_reg_3_ ( .J(n84), .K(n84), .TI(N116), .TE(N115), .CP(clk), .Q(hh[7]), .QN(n6) );
  GTECH_FJK1S hh_ones_reg_0_ ( .J(n84), .K(n84), .TI(N88), .TE(N91), .CP(clk), 
        .Q(hh[0]), .QN(n7) );
  GTECH_FJK1S hh_ones_reg_1_ ( .J(n84), .K(n84), .TI(N89), .TE(N91), .CP(clk), 
        .Q(hh[1]), .QN(n109) );
  GTECH_FJK1S hh_ones_reg_2_ ( .J(n84), .K(n84), .TI(N90), .TE(N91), .CP(clk), 
        .Q(hh[2]), .QN(n125) );
  GTECH_FJK1S hh_ones_reg_3_ ( .J(n84), .K(n84), .TI(N92), .TE(N91), .CP(clk), 
        .Q(hh[3]), .QN(n124) );
  GTECH_FJK1S hh_tens_reg_1_ ( .J(n84), .K(n84), .TI(N112), .TE(N115), .CP(clk), .Q(hh[5]), .QN(n8) );
  GTECH_FJK1S pm_temp_reg ( .J(n84), .K(n84), .TI(N122), .TE(N121), .CP(clk), 
        .Q(pm), .QN(n9) );
  GTECH_ZERO U134 ( .Z(n84) );
  GTECH_AND2 U135 ( .A(n126), .B(n127), .Z(N92) );
  GTECH_XOR2 U136 ( .A(n128), .B(n124), .Z(n126) );
  GTECH_OR_NOT U137 ( .A(n129), .B(n130), .Z(n128) );
  GTECH_NAND2 U138 ( .A(n131), .B(n132), .Z(N91) );
  GTECH_AND2 U139 ( .A(n133), .B(n127), .Z(N90) );
  GTECH_NOT U140 ( .A(n134), .Z(n127) );
  GTECH_XOR2 U141 ( .A(n129), .B(n125), .Z(n133) );
  GTECH_NAND2 U142 ( .A(n135), .B(n136), .Z(n129) );
  GTECH_OAI21 U143 ( .A(n137), .B(n134), .C(n131), .Z(N89) );
  GTECH_XOR2 U144 ( .A(n136), .B(n7), .Z(n137) );
  GTECH_OAI22 U145 ( .A(n132), .B(n138), .C(n135), .D(n134), .Z(N88) );
  GTECH_NAND3 U146 ( .A(n138), .B(n139), .C(n140), .Z(n134) );
  GTECH_MUX2 U147 ( .A(n141), .B(n142), .S(n110), .Z(N75) );
  GTECH_AND2 U148 ( .A(n143), .B(n144), .Z(n142) );
  GTECH_OAI21 U149 ( .A(n145), .B(n144), .C(n146), .Z(n141) );
  GTECH_NOT U150 ( .A(n147), .Z(n146) );
  GTECH_NOT U151 ( .A(n111), .Z(n144) );
  GTECH_MUX2 U152 ( .A(n147), .B(n148), .S(n111), .Z(N73) );
  GTECH_AND2 U153 ( .A(n143), .B(n149), .Z(n148) );
  GTECH_OAI21 U154 ( .A(n149), .B(n145), .C(n150), .Z(n147) );
  GTECH_MUX2 U155 ( .A(N71), .B(n143), .S(n112), .Z(N72) );
  GTECH_NOT U156 ( .A(n151), .Z(n143) );
  GTECH_NAND2 U157 ( .A(n152), .B(n153), .Z(n151) );
  GTECH_NOT U158 ( .A(n3), .Z(n153) );
  GTECH_NOT U159 ( .A(n150), .Z(N71) );
  GTECH_NAND2 U160 ( .A(n3), .B(n152), .Z(n150) );
  GTECH_NOT U161 ( .A(n145), .Z(n152) );
  GTECH_NAND3 U162 ( .A(n154), .B(n131), .C(n155), .Z(n145) );
  GTECH_NOT U163 ( .A(n156), .Z(n155) );
  GTECH_MUX2 U164 ( .A(n157), .B(n158), .S(n113), .Z(N59) );
  GTECH_AND2 U165 ( .A(n159), .B(n160), .Z(n158) );
  GTECH_OAI21 U166 ( .A(n160), .B(n161), .C(n162), .Z(n157) );
  GTECH_NOT U167 ( .A(n163), .Z(n162) );
  GTECH_MUX2 U168 ( .A(n163), .B(n159), .S(n116), .Z(N57) );
  GTECH_NOT U169 ( .A(n164), .Z(n159) );
  GTECH_NAND3 U170 ( .A(n165), .B(n166), .C(n167), .Z(n164) );
  GTECH_OAI21 U171 ( .A(n166), .B(n161), .C(n168), .Z(n163) );
  GTECH_MUX2 U172 ( .A(N55), .B(n169), .S(n115), .Z(N56) );
  GTECH_AND2 U173 ( .A(n167), .B(n165), .Z(n169) );
  GTECH_NOT U174 ( .A(n114), .Z(n165) );
  GTECH_NOT U175 ( .A(n168), .Z(N55) );
  GTECH_NAND2 U176 ( .A(n114), .B(n167), .Z(n168) );
  GTECH_NOT U177 ( .A(n161), .Z(n167) );
  GTECH_NAND2 U178 ( .A(n170), .B(n171), .Z(n161) );
  GTECH_NOT U179 ( .A(N74), .Z(n171) );
  GTECH_NAND2 U180 ( .A(n131), .B(n156), .Z(N74) );
  GTECH_NOT U181 ( .A(n172), .Z(n170) );
  GTECH_MUX2 U182 ( .A(n173), .B(n174), .S(ss[7]), .Z(N43) );
  GTECH_OAI21 U183 ( .A(ss[6]), .B(n175), .C(n176), .Z(n174) );
  GTECH_NOT U184 ( .A(n177), .Z(n176) );
  GTECH_AND2 U185 ( .A(n178), .B(ss[6]), .Z(n173) );
  GTECH_MUX2 U186 ( .A(n179), .B(n177), .S(ss[6]), .Z(N41) );
  GTECH_OAI21 U187 ( .A(ss[5]), .B(n175), .C(n180), .Z(n177) );
  GTECH_AND2 U188 ( .A(ss[5]), .B(n178), .Z(n179) );
  GTECH_MUX2 U189 ( .A(n178), .B(N39), .S(ss[5]), .Z(N40) );
  GTECH_NOT U190 ( .A(n181), .Z(n178) );
  GTECH_NAND2 U191 ( .A(n182), .B(ss[4]), .Z(n181) );
  GTECH_NOT U192 ( .A(n180), .Z(N39) );
  GTECH_NAND2 U193 ( .A(n182), .B(n183), .Z(n180) );
  GTECH_NOT U194 ( .A(n175), .Z(n182) );
  GTECH_NAND2 U195 ( .A(n184), .B(n185), .Z(n175) );
  GTECH_NOT U196 ( .A(N58), .Z(n185) );
  GTECH_NAND2 U197 ( .A(n131), .B(n172), .Z(N58) );
  GTECH_NOT U198 ( .A(n186), .Z(n184) );
  GTECH_MUX2 U199 ( .A(n187), .B(n188), .S(ss[3]), .Z(N26) );
  GTECH_OAI21 U200 ( .A(ss[2]), .B(n189), .C(n190), .Z(n188) );
  GTECH_NOT U201 ( .A(n191), .Z(n190) );
  GTECH_AND2 U202 ( .A(ss[2]), .B(n192), .Z(n187) );
  GTECH_NAND2 U203 ( .A(n131), .B(n193), .Z(N25) );
  GTECH_MUX2 U204 ( .A(n192), .B(n191), .S(ss[2]), .Z(N24) );
  GTECH_OAI21 U205 ( .A(ss[1]), .B(n189), .C(n194), .Z(n191) );
  GTECH_NOT U206 ( .A(n195), .Z(n192) );
  GTECH_NAND3 U207 ( .A(n196), .B(ss[0]), .C(ss[1]), .Z(n195) );
  GTECH_MUX2 U208 ( .A(n197), .B(N22), .S(ss[1]), .Z(N23) );
  GTECH_AND2 U209 ( .A(n196), .B(ss[0]), .Z(n197) );
  GTECH_NOT U210 ( .A(n194), .Z(N22) );
  GTECH_NAND2 U211 ( .A(n196), .B(n198), .Z(n194) );
  GTECH_NOT U212 ( .A(n189), .Z(n196) );
  GTECH_NAND2 U213 ( .A(ena), .B(n199), .Z(n189) );
  GTECH_NOT U214 ( .A(N42), .Z(n199) );
  GTECH_NAND2 U215 ( .A(n131), .B(n186), .Z(N42) );
  GTECH_AND2 U216 ( .A(n200), .B(n9), .Z(N122) );
  GTECH_NOT U217 ( .A(n201), .Z(n200) );
  GTECH_NAND2 U218 ( .A(n131), .B(n201), .Z(N121) );
  GTECH_NAND4 U219 ( .A(n140), .B(n202), .C(n109), .D(n135), .Z(n201) );
  GTECH_NOT U220 ( .A(n7), .Z(n135) );
  GTECH_AND2 U221 ( .A(n203), .B(n204), .Z(N116) );
  GTECH_XOR2 U222 ( .A(n205), .B(n6), .Z(n203) );
  GTECH_OR2 U223 ( .A(n5), .B(n206), .Z(n205) );
  GTECH_NAND3 U224 ( .A(n139), .B(n131), .C(n138), .Z(N115) );
  GTECH_NAND4 U225 ( .A(n7), .B(n202), .C(n207), .D(n136), .Z(n138) );
  GTECH_AND3 U226 ( .A(n6), .B(n5), .C(n208), .Z(n202) );
  GTECH_AND4 U227 ( .A(n209), .B(n124), .C(n125), .D(n8), .Z(n208) );
  GTECH_AND2 U228 ( .A(n210), .B(n204), .Z(N114) );
  GTECH_XOR2 U229 ( .A(n206), .B(n5), .Z(n210) );
  GTECH_NAND2 U230 ( .A(n211), .B(n209), .Z(n206) );
  GTECH_NOT U231 ( .A(n8), .Z(n211) );
  GTECH_AND2 U232 ( .A(n204), .B(n212), .Z(N112) );
  GTECH_XOR2 U233 ( .A(n8), .B(n4), .Z(n212) );
  GTECH_NOT U234 ( .A(n213), .Z(n204) );
  GTECH_OAI21 U235 ( .A(n213), .B(n209), .C(n131), .Z(N110) );
  GTECH_NOT U236 ( .A(n4), .Z(n209) );
  GTECH_NAND2 U237 ( .A(n214), .B(n140), .Z(n213) );
  GTECH_NOT U238 ( .A(n132), .Z(n140) );
  GTECH_NAND2 U239 ( .A(n207), .B(n131), .Z(n132) );
  GTECH_NOT U240 ( .A(reset), .Z(n131) );
  GTECH_NOT U241 ( .A(n154), .Z(n207) );
  GTECH_NOT U242 ( .A(n139), .Z(n214) );
  GTECH_OR5 U243 ( .A(n7), .B(n124), .C(n154), .D(n136), .E(n130), .Z(n139) );
  GTECH_NOT U244 ( .A(n125), .Z(n130) );
  GTECH_NOT U245 ( .A(n109), .Z(n136) );
  GTECH_OR5 U246 ( .A(n3), .B(n111), .C(n156), .D(n215), .E(n149), .Z(n154) );
  GTECH_NOT U247 ( .A(n112), .Z(n149) );
  GTECH_NOT U248 ( .A(n110), .Z(n215) );
  GTECH_OR5 U249 ( .A(n114), .B(n113), .C(n172), .D(n166), .E(n160), .Z(n156)
         );
  GTECH_NOT U250 ( .A(n116), .Z(n160) );
  GTECH_NOT U251 ( .A(n115), .Z(n166) );
  GTECH_OR5 U252 ( .A(ss[7]), .B(ss[5]), .C(n186), .D(n183), .E(n216), .Z(n172) );
  GTECH_NOT U253 ( .A(ss[6]), .Z(n216) );
  GTECH_NOT U254 ( .A(ss[4]), .Z(n183) );
  GTECH_OR5 U255 ( .A(ss[2]), .B(ss[1]), .C(n193), .D(n198), .E(n217), .Z(n186) );
  GTECH_NOT U256 ( .A(ss[3]), .Z(n217) );
  GTECH_NOT U257 ( .A(ss[0]), .Z(n198) );
  GTECH_NOT U258 ( .A(ena), .Z(n193) );
endmodule

