
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI2N2 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_OR_NOT U83 ( .A(n97), .B(n93), .Z(n96) );
  GTECH_XOR2 U84 ( .A(n90), .B(n98), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n98) );
  GTECH_OAI21 U86 ( .A(n99), .B(n100), .C(n101), .Z(n89) );
  GTECH_OAI21 U87 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  GTECH_OR_NOT U88 ( .A(n105), .B(I_b[7]), .Z(n90) );
  GTECH_NOT U89 ( .A(n106), .Z(n84) );
  GTECH_OR_NOT U90 ( .A(n107), .B(n108), .Z(n106) );
  GTECH_XOR2 U91 ( .A(n109), .B(n108), .Z(N153) );
  GTECH_NOT U92 ( .A(n110), .Z(n108) );
  GTECH_XNOR3 U93 ( .A(n97), .B(n93), .C(n111), .Z(n110) );
  GTECH_NOT U94 ( .A(n95), .Z(n111) );
  GTECH_XNOR3 U95 ( .A(n102), .B(n104), .C(n99), .Z(n95) );
  GTECH_NOT U96 ( .A(n103), .Z(n99) );
  GTECH_OAI21 U97 ( .A(n112), .B(n113), .C(n114), .Z(n103) );
  GTECH_OAI21 U98 ( .A(n115), .B(n116), .C(n117), .Z(n114) );
  GTECH_NOT U99 ( .A(n118), .Z(n104) );
  GTECH_OR_NOT U100 ( .A(n119), .B(I_b[7]), .Z(n118) );
  GTECH_NOT U101 ( .A(n100), .Z(n102) );
  GTECH_OR_NOT U102 ( .A(n120), .B(I_a[7]), .Z(n100) );
  GTECH_NOT U103 ( .A(I_b[6]), .Z(n120) );
  GTECH_ADD_ABC U104 ( .A(n121), .B(n122), .C(n123), .COUT(n93) );
  GTECH_NOT U105 ( .A(n124), .Z(n123) );
  GTECH_XOR2 U106 ( .A(n125), .B(n126), .Z(n122) );
  GTECH_AND2 U107 ( .A(I_a[7]), .B(I_b[5]), .Z(n126) );
  GTECH_NOT U108 ( .A(n94), .Z(n97) );
  GTECH_OR_NOT U109 ( .A(n125), .B(I_a[7]), .Z(n94) );
  GTECH_NOT U110 ( .A(n107), .Z(n109) );
  GTECH_OR_NOT U111 ( .A(n127), .B(n128), .Z(n107) );
  GTECH_XOR2 U112 ( .A(n127), .B(n129), .Z(N152) );
  GTECH_NOT U113 ( .A(n128), .Z(n129) );
  GTECH_XOR4 U114 ( .A(n130), .B(n125), .C(n124), .D(n121), .Z(n128) );
  GTECH_ADD_ABC U115 ( .A(n131), .B(n132), .C(n133), .COUT(n121) );
  GTECH_XNOR3 U116 ( .A(n134), .B(n135), .C(n136), .Z(n132) );
  GTECH_XNOR3 U117 ( .A(n115), .B(n117), .C(n112), .Z(n124) );
  GTECH_NOT U118 ( .A(n116), .Z(n112) );
  GTECH_OAI21 U119 ( .A(n137), .B(n138), .C(n139), .Z(n116) );
  GTECH_OAI21 U120 ( .A(n140), .B(n141), .C(n142), .Z(n139) );
  GTECH_NOT U121 ( .A(n143), .Z(n117) );
  GTECH_OR_NOT U122 ( .A(n144), .B(I_b[7]), .Z(n143) );
  GTECH_NOT U123 ( .A(n113), .Z(n115) );
  GTECH_OR_NOT U124 ( .A(n119), .B(I_b[6]), .Z(n113) );
  GTECH_NOT U125 ( .A(I_a[6]), .Z(n119) );
  GTECH_OA21 U126 ( .A(n145), .B(n146), .C(n147), .Z(n125) );
  GTECH_OAI21 U127 ( .A(n134), .B(n136), .C(n135), .Z(n147) );
  GTECH_AND2 U128 ( .A(I_b[5]), .B(I_a[7]), .Z(n130) );
  GTECH_ADD_ABC U129 ( .A(n148), .B(n149), .C(n150), .COUT(n127) );
  GTECH_OA22 U130 ( .A(n151), .B(n105), .C(n152), .D(n153), .Z(n149) );
  GTECH_OA21 U131 ( .A(n154), .B(n155), .C(n156), .Z(n148) );
  GTECH_XNOR3 U132 ( .A(n157), .B(n150), .C(n158), .Z(N151) );
  GTECH_OA21 U133 ( .A(n154), .B(n155), .C(n156), .Z(n158) );
  GTECH_OAI21 U134 ( .A(n159), .B(n160), .C(n161), .Z(n156) );
  GTECH_XOR2 U135 ( .A(n131), .B(n162), .Z(n150) );
  GTECH_XOR4 U136 ( .A(n135), .B(n145), .C(n133), .D(n134), .Z(n162) );
  GTECH_NOT U137 ( .A(n146), .Z(n134) );
  GTECH_OR_NOT U138 ( .A(n163), .B(I_a[7]), .Z(n146) );
  GTECH_NOT U139 ( .A(n164), .Z(n133) );
  GTECH_XNOR3 U140 ( .A(n140), .B(n142), .C(n137), .Z(n164) );
  GTECH_NOT U141 ( .A(n141), .Z(n137) );
  GTECH_OAI21 U142 ( .A(n165), .B(n166), .C(n167), .Z(n141) );
  GTECH_OAI21 U143 ( .A(n168), .B(n169), .C(n170), .Z(n167) );
  GTECH_NOT U144 ( .A(n171), .Z(n142) );
  GTECH_OR_NOT U145 ( .A(n172), .B(I_b[7]), .Z(n171) );
  GTECH_NOT U146 ( .A(n138), .Z(n140) );
  GTECH_OR_NOT U147 ( .A(n144), .B(I_b[6]), .Z(n138) );
  GTECH_NOT U148 ( .A(I_a[5]), .Z(n144) );
  GTECH_NOT U149 ( .A(n136), .Z(n145) );
  GTECH_OAI21 U150 ( .A(n173), .B(n174), .C(n175), .Z(n136) );
  GTECH_OAI21 U151 ( .A(n176), .B(n177), .C(n178), .Z(n175) );
  GTECH_NOT U152 ( .A(n179), .Z(n135) );
  GTECH_OR_NOT U153 ( .A(n180), .B(I_a[6]), .Z(n179) );
  GTECH_ADD_ABC U154 ( .A(n181), .B(n182), .C(n183), .COUT(n131) );
  GTECH_NOT U155 ( .A(n184), .Z(n183) );
  GTECH_XNOR3 U156 ( .A(n176), .B(n178), .C(n177), .Z(n182) );
  GTECH_OA22 U157 ( .A(n151), .B(n105), .C(n152), .D(n153), .Z(n157) );
  GTECH_NOT U158 ( .A(n185), .Z(n153) );
  GTECH_NOT U159 ( .A(I_a[7]), .Z(n105) );
  GTECH_XNOR3 U160 ( .A(n154), .B(n159), .C(n161), .Z(N150) );
  GTECH_XOR2 U161 ( .A(n186), .B(n181), .Z(n161) );
  GTECH_ADD_ABC U162 ( .A(n187), .B(n188), .C(n189), .COUT(n181) );
  GTECH_NOT U163 ( .A(n190), .Z(n189) );
  GTECH_XNOR3 U164 ( .A(n191), .B(n192), .C(n193), .Z(n188) );
  GTECH_XOR4 U165 ( .A(n178), .B(n173), .C(n184), .D(n176), .Z(n186) );
  GTECH_NOT U166 ( .A(n174), .Z(n176) );
  GTECH_OR_NOT U167 ( .A(n163), .B(I_a[6]), .Z(n174) );
  GTECH_XNOR3 U168 ( .A(n168), .B(n170), .C(n165), .Z(n184) );
  GTECH_NOT U169 ( .A(n169), .Z(n165) );
  GTECH_OAI21 U170 ( .A(n194), .B(n195), .C(n196), .Z(n169) );
  GTECH_OAI21 U171 ( .A(n197), .B(n198), .C(n199), .Z(n196) );
  GTECH_NOT U172 ( .A(n200), .Z(n170) );
  GTECH_OR_NOT U173 ( .A(n201), .B(I_b[7]), .Z(n200) );
  GTECH_NOT U174 ( .A(n166), .Z(n168) );
  GTECH_OR_NOT U175 ( .A(n172), .B(I_b[6]), .Z(n166) );
  GTECH_NOT U176 ( .A(n177), .Z(n173) );
  GTECH_OAI21 U177 ( .A(n202), .B(n203), .C(n204), .Z(n177) );
  GTECH_OAI21 U178 ( .A(n191), .B(n193), .C(n192), .Z(n204) );
  GTECH_NOT U179 ( .A(n205), .Z(n178) );
  GTECH_OR_NOT U180 ( .A(n180), .B(I_a[5]), .Z(n205) );
  GTECH_NOT U181 ( .A(I_b[5]), .Z(n180) );
  GTECH_NOT U182 ( .A(n155), .Z(n159) );
  GTECH_XOR2 U183 ( .A(n185), .B(n152), .Z(n155) );
  GTECH_AOI2N2 U184 ( .A(n206), .B(n207), .C(n208), .D(n209), .Z(n152) );
  GTECH_OR_NOT U185 ( .A(n210), .B(n208), .Z(n207) );
  GTECH_XOR2 U186 ( .A(n211), .B(n151), .Z(n185) );
  GTECH_OA21 U187 ( .A(n212), .B(n213), .C(n214), .Z(n151) );
  GTECH_OAI21 U188 ( .A(n215), .B(n216), .C(n217), .Z(n214) );
  GTECH_OR_NOT U189 ( .A(n218), .B(I_a[7]), .Z(n211) );
  GTECH_NOT U190 ( .A(n160), .Z(n154) );
  GTECH_OAI2N2 U191 ( .A(n219), .B(n220), .C(n221), .D(n222), .Z(n160) );
  GTECH_OR_NOT U192 ( .A(n223), .B(n219), .Z(n222) );
  GTECH_XNOR3 U193 ( .A(n219), .B(n223), .C(n221), .Z(N149) );
  GTECH_XOR2 U194 ( .A(n224), .B(n187), .Z(n221) );
  GTECH_ADD_ABC U195 ( .A(n225), .B(n226), .C(n227), .COUT(n187) );
  GTECH_XNOR3 U196 ( .A(n228), .B(n229), .C(n230), .Z(n226) );
  GTECH_OA21 U197 ( .A(n231), .B(n232), .C(n233), .Z(n225) );
  GTECH_XOR4 U198 ( .A(n192), .B(n202), .C(n190), .D(n191), .Z(n224) );
  GTECH_NOT U199 ( .A(n203), .Z(n191) );
  GTECH_OR_NOT U200 ( .A(n163), .B(I_a[5]), .Z(n203) );
  GTECH_NOT U201 ( .A(I_b[4]), .Z(n163) );
  GTECH_XNOR3 U202 ( .A(n197), .B(n199), .C(n194), .Z(n190) );
  GTECH_NOT U203 ( .A(n198), .Z(n194) );
  GTECH_OAI21 U204 ( .A(n234), .B(n235), .C(n236), .Z(n198) );
  GTECH_NOT U205 ( .A(n237), .Z(n199) );
  GTECH_OR_NOT U206 ( .A(n238), .B(I_b[7]), .Z(n237) );
  GTECH_NOT U207 ( .A(n195), .Z(n197) );
  GTECH_OR_NOT U208 ( .A(n201), .B(I_b[6]), .Z(n195) );
  GTECH_NOT U209 ( .A(n193), .Z(n202) );
  GTECH_OAI21 U210 ( .A(n239), .B(n240), .C(n241), .Z(n193) );
  GTECH_OAI21 U211 ( .A(n228), .B(n230), .C(n229), .Z(n241) );
  GTECH_NOT U212 ( .A(n242), .Z(n192) );
  GTECH_OR_NOT U213 ( .A(n172), .B(I_b[5]), .Z(n242) );
  GTECH_NOT U214 ( .A(n220), .Z(n223) );
  GTECH_XNOR3 U215 ( .A(n210), .B(n208), .C(n243), .Z(n220) );
  GTECH_NOT U216 ( .A(n206), .Z(n243) );
  GTECH_XNOR3 U217 ( .A(n215), .B(n217), .C(n212), .Z(n206) );
  GTECH_NOT U218 ( .A(n216), .Z(n212) );
  GTECH_OAI21 U219 ( .A(n244), .B(n245), .C(n246), .Z(n216) );
  GTECH_OAI21 U220 ( .A(n247), .B(n248), .C(n249), .Z(n246) );
  GTECH_NOT U221 ( .A(n250), .Z(n217) );
  GTECH_OR_NOT U222 ( .A(n218), .B(I_a[6]), .Z(n250) );
  GTECH_NOT U223 ( .A(n213), .Z(n215) );
  GTECH_OR_NOT U224 ( .A(n251), .B(I_a[7]), .Z(n213) );
  GTECH_ADD_ABC U225 ( .A(n252), .B(n253), .C(n254), .COUT(n208) );
  GTECH_NOT U226 ( .A(n255), .Z(n254) );
  GTECH_XOR2 U227 ( .A(n256), .B(n257), .Z(n253) );
  GTECH_AND2 U228 ( .A(I_a[7]), .B(I_b[1]), .Z(n257) );
  GTECH_NOT U229 ( .A(n209), .Z(n210) );
  GTECH_OR_NOT U230 ( .A(n256), .B(I_a[7]), .Z(n209) );
  GTECH_ADD_ABC U231 ( .A(n258), .B(n259), .C(n260), .COUT(n219) );
  GTECH_XNOR3 U232 ( .A(n252), .B(n261), .C(n255), .Z(n259) );
  GTECH_XOR2 U233 ( .A(n262), .B(n258), .Z(N148) );
  GTECH_ADD_ABC U234 ( .A(n263), .B(n264), .C(n265), .COUT(n258) );
  GTECH_NOT U235 ( .A(n266), .Z(n265) );
  GTECH_XNOR3 U236 ( .A(n267), .B(n268), .C(n269), .Z(n264) );
  GTECH_XOR4 U237 ( .A(n261), .B(n252), .C(n255), .D(n260), .Z(n262) );
  GTECH_XOR2 U238 ( .A(n270), .B(n271), .Z(n260) );
  GTECH_XOR4 U239 ( .A(n229), .B(n239), .C(n227), .D(n228), .Z(n271) );
  GTECH_NOT U240 ( .A(n240), .Z(n228) );
  GTECH_OR_NOT U241 ( .A(n172), .B(I_b[4]), .Z(n240) );
  GTECH_XNOR3 U242 ( .A(n272), .B(n273), .C(n274), .Z(n227) );
  GTECH_NOT U243 ( .A(n236), .Z(n274) );
  GTECH_NAND3 U244 ( .A(I_b[6]), .B(I_a[1]), .C(n275), .Z(n236) );
  GTECH_NOT U245 ( .A(n235), .Z(n273) );
  GTECH_OR_NOT U246 ( .A(n276), .B(I_b[7]), .Z(n235) );
  GTECH_NOT U247 ( .A(n234), .Z(n272) );
  GTECH_OR_NOT U248 ( .A(n238), .B(I_b[6]), .Z(n234) );
  GTECH_NOT U249 ( .A(n230), .Z(n239) );
  GTECH_OAI21 U250 ( .A(n277), .B(n278), .C(n279), .Z(n230) );
  GTECH_OAI21 U251 ( .A(n280), .B(n281), .C(n282), .Z(n279) );
  GTECH_NOT U252 ( .A(n283), .Z(n229) );
  GTECH_OR_NOT U253 ( .A(n201), .B(I_b[5]), .Z(n283) );
  GTECH_OA21 U254 ( .A(n231), .B(n232), .C(n233), .Z(n270) );
  GTECH_OAI21 U255 ( .A(n284), .B(n285), .C(n286), .Z(n233) );
  GTECH_XNOR3 U256 ( .A(n247), .B(n249), .C(n244), .Z(n255) );
  GTECH_NOT U257 ( .A(n248), .Z(n244) );
  GTECH_OAI21 U258 ( .A(n287), .B(n288), .C(n289), .Z(n248) );
  GTECH_OAI21 U259 ( .A(n290), .B(n291), .C(n292), .Z(n289) );
  GTECH_NOT U260 ( .A(n293), .Z(n249) );
  GTECH_OR_NOT U261 ( .A(n218), .B(I_a[5]), .Z(n293) );
  GTECH_NOT U262 ( .A(I_b[3]), .Z(n218) );
  GTECH_NOT U263 ( .A(n245), .Z(n247) );
  GTECH_OR_NOT U264 ( .A(n251), .B(I_a[6]), .Z(n245) );
  GTECH_ADD_ABC U265 ( .A(n267), .B(n294), .C(n295), .COUT(n252) );
  GTECH_XNOR3 U266 ( .A(n296), .B(n297), .C(n298), .Z(n294) );
  GTECH_XOR2 U267 ( .A(n299), .B(n256), .Z(n261) );
  GTECH_OA21 U268 ( .A(n300), .B(n301), .C(n302), .Z(n256) );
  GTECH_OAI21 U269 ( .A(n296), .B(n298), .C(n297), .Z(n302) );
  GTECH_AND2 U270 ( .A(I_b[1]), .B(I_a[7]), .Z(n299) );
  GTECH_XOR2 U271 ( .A(n303), .B(n263), .Z(N147) );
  GTECH_ADD_ABC U272 ( .A(n304), .B(n305), .C(n306), .COUT(n263) );
  GTECH_XNOR3 U273 ( .A(n307), .B(n308), .C(n309), .Z(n305) );
  GTECH_OA21 U274 ( .A(n310), .B(n311), .C(n312), .Z(n304) );
  GTECH_XOR4 U275 ( .A(n268), .B(n295), .C(n266), .D(n267), .Z(n303) );
  GTECH_ADD_ABC U276 ( .A(n307), .B(n313), .C(n314), .COUT(n267) );
  GTECH_NOT U277 ( .A(n309), .Z(n314) );
  GTECH_XNOR3 U278 ( .A(n315), .B(n316), .C(n317), .Z(n313) );
  GTECH_XNOR3 U279 ( .A(n286), .B(n232), .C(n285), .Z(n266) );
  GTECH_NOT U280 ( .A(n231), .Z(n285) );
  GTECH_XOR2 U281 ( .A(n318), .B(n275), .Z(n231) );
  GTECH_NOT U282 ( .A(n319), .Z(n275) );
  GTECH_OR_NOT U283 ( .A(n320), .B(I_b[7]), .Z(n319) );
  GTECH_OR_NOT U284 ( .A(n276), .B(I_b[6]), .Z(n318) );
  GTECH_NOT U285 ( .A(n284), .Z(n232) );
  GTECH_XNOR3 U286 ( .A(n280), .B(n282), .C(n277), .Z(n284) );
  GTECH_NOT U287 ( .A(n281), .Z(n277) );
  GTECH_OAI21 U288 ( .A(n321), .B(n322), .C(n323), .Z(n281) );
  GTECH_NOT U289 ( .A(n324), .Z(n282) );
  GTECH_OR_NOT U290 ( .A(n238), .B(I_b[5]), .Z(n324) );
  GTECH_NOT U291 ( .A(n278), .Z(n280) );
  GTECH_OR_NOT U292 ( .A(n201), .B(I_b[4]), .Z(n278) );
  GTECH_NOT U293 ( .A(n325), .Z(n286) );
  GTECH_NAND3 U294 ( .A(I_a[0]), .B(n326), .C(I_b[6]), .Z(n325) );
  GTECH_NOT U295 ( .A(n327), .Z(n326) );
  GTECH_NOT U296 ( .A(n269), .Z(n295) );
  GTECH_XNOR3 U297 ( .A(n290), .B(n292), .C(n287), .Z(n269) );
  GTECH_NOT U298 ( .A(n291), .Z(n287) );
  GTECH_OAI21 U299 ( .A(n328), .B(n329), .C(n330), .Z(n291) );
  GTECH_OAI21 U300 ( .A(n331), .B(n332), .C(n333), .Z(n330) );
  GTECH_NOT U301 ( .A(n334), .Z(n292) );
  GTECH_OR_NOT U302 ( .A(n172), .B(I_b[3]), .Z(n334) );
  GTECH_NOT U303 ( .A(n288), .Z(n290) );
  GTECH_OR_NOT U304 ( .A(n251), .B(I_a[5]), .Z(n288) );
  GTECH_NOT U305 ( .A(I_b[2]), .Z(n251) );
  GTECH_NOT U306 ( .A(n335), .Z(n268) );
  GTECH_XNOR3 U307 ( .A(n296), .B(n297), .C(n300), .Z(n335) );
  GTECH_NOT U308 ( .A(n298), .Z(n300) );
  GTECH_OAI21 U309 ( .A(n336), .B(n337), .C(n338), .Z(n298) );
  GTECH_OAI21 U310 ( .A(n315), .B(n317), .C(n316), .Z(n338) );
  GTECH_NOT U311 ( .A(n339), .Z(n297) );
  GTECH_OR_NOT U312 ( .A(n340), .B(I_a[6]), .Z(n339) );
  GTECH_NOT U313 ( .A(n301), .Z(n296) );
  GTECH_OR_NOT U314 ( .A(n341), .B(I_a[7]), .Z(n301) );
  GTECH_XOR2 U315 ( .A(n342), .B(n343), .Z(N146) );
  GTECH_OA21 U316 ( .A(n310), .B(n311), .C(n312), .Z(n343) );
  GTECH_OAI21 U317 ( .A(n344), .B(n345), .C(n346), .Z(n312) );
  GTECH_XOR4 U318 ( .A(n308), .B(n307), .C(n309), .D(n306), .Z(n342) );
  GTECH_XOR2 U319 ( .A(n327), .B(n347), .Z(n306) );
  GTECH_AND2 U320 ( .A(I_b[6]), .B(I_a[0]), .Z(n347) );
  GTECH_XNOR3 U321 ( .A(n348), .B(n349), .C(n350), .Z(n327) );
  GTECH_NOT U322 ( .A(n323), .Z(n350) );
  GTECH_NAND3 U323 ( .A(I_b[4]), .B(I_a[1]), .C(n351), .Z(n323) );
  GTECH_NOT U324 ( .A(n322), .Z(n349) );
  GTECH_OR_NOT U325 ( .A(n276), .B(I_b[5]), .Z(n322) );
  GTECH_NOT U326 ( .A(n321), .Z(n348) );
  GTECH_OR_NOT U327 ( .A(n238), .B(I_b[4]), .Z(n321) );
  GTECH_XNOR3 U328 ( .A(n331), .B(n333), .C(n328), .Z(n309) );
  GTECH_NOT U329 ( .A(n332), .Z(n328) );
  GTECH_OAI21 U330 ( .A(n352), .B(n353), .C(n354), .Z(n332) );
  GTECH_OAI21 U331 ( .A(n355), .B(n356), .C(n357), .Z(n354) );
  GTECH_NOT U332 ( .A(n358), .Z(n333) );
  GTECH_OR_NOT U333 ( .A(n201), .B(I_b[3]), .Z(n358) );
  GTECH_NOT U334 ( .A(n329), .Z(n331) );
  GTECH_OR_NOT U335 ( .A(n172), .B(I_b[2]), .Z(n329) );
  GTECH_NOT U336 ( .A(I_a[4]), .Z(n172) );
  GTECH_ADD_ABC U337 ( .A(n359), .B(n360), .C(n361), .COUT(n307) );
  GTECH_NOT U338 ( .A(n362), .Z(n361) );
  GTECH_XNOR3 U339 ( .A(n363), .B(n364), .C(n365), .Z(n360) );
  GTECH_NOT U340 ( .A(n366), .Z(n308) );
  GTECH_XNOR3 U341 ( .A(n315), .B(n316), .C(n336), .Z(n366) );
  GTECH_NOT U342 ( .A(n317), .Z(n336) );
  GTECH_OAI21 U343 ( .A(n367), .B(n368), .C(n369), .Z(n317) );
  GTECH_OAI21 U344 ( .A(n363), .B(n365), .C(n364), .Z(n369) );
  GTECH_NOT U345 ( .A(n370), .Z(n316) );
  GTECH_OR_NOT U346 ( .A(n340), .B(I_a[5]), .Z(n370) );
  GTECH_NOT U347 ( .A(n337), .Z(n315) );
  GTECH_OR_NOT U348 ( .A(n341), .B(I_a[6]), .Z(n337) );
  GTECH_XNOR3 U349 ( .A(n346), .B(n311), .C(n345), .Z(N145) );
  GTECH_NOT U350 ( .A(n310), .Z(n345) );
  GTECH_XOR2 U351 ( .A(n371), .B(n351), .Z(n310) );
  GTECH_NOT U352 ( .A(n372), .Z(n351) );
  GTECH_OR_NOT U353 ( .A(n320), .B(I_b[5]), .Z(n372) );
  GTECH_OR_NOT U354 ( .A(n276), .B(I_b[4]), .Z(n371) );
  GTECH_NOT U355 ( .A(n344), .Z(n311) );
  GTECH_XOR2 U356 ( .A(n373), .B(n359), .Z(n344) );
  GTECH_ADD_ABC U357 ( .A(n374), .B(n375), .C(n376), .COUT(n359) );
  GTECH_XNOR3 U358 ( .A(n377), .B(n378), .C(n379), .Z(n375) );
  GTECH_OA21 U359 ( .A(n380), .B(n381), .C(n382), .Z(n374) );
  GTECH_XOR4 U360 ( .A(n364), .B(n367), .C(n362), .D(n363), .Z(n373) );
  GTECH_NOT U361 ( .A(n368), .Z(n363) );
  GTECH_OR_NOT U362 ( .A(n341), .B(I_a[5]), .Z(n368) );
  GTECH_XNOR3 U363 ( .A(n355), .B(n357), .C(n352), .Z(n362) );
  GTECH_NOT U364 ( .A(n356), .Z(n352) );
  GTECH_OAI21 U365 ( .A(n383), .B(n384), .C(n385), .Z(n356) );
  GTECH_NOT U366 ( .A(n386), .Z(n357) );
  GTECH_OR_NOT U367 ( .A(n238), .B(I_b[3]), .Z(n386) );
  GTECH_NOT U368 ( .A(n353), .Z(n355) );
  GTECH_OR_NOT U369 ( .A(n201), .B(I_b[2]), .Z(n353) );
  GTECH_NOT U370 ( .A(n365), .Z(n367) );
  GTECH_OAI21 U371 ( .A(n387), .B(n388), .C(n389), .Z(n365) );
  GTECH_OAI21 U372 ( .A(n377), .B(n379), .C(n378), .Z(n389) );
  GTECH_NOT U373 ( .A(n388), .Z(n377) );
  GTECH_NOT U374 ( .A(n390), .Z(n364) );
  GTECH_OR_NOT U375 ( .A(n340), .B(I_a[4]), .Z(n390) );
  GTECH_NOT U376 ( .A(n391), .Z(n346) );
  GTECH_NAND3 U377 ( .A(I_a[0]), .B(n392), .C(I_b[4]), .Z(n391) );
  GTECH_XOR2 U378 ( .A(n393), .B(n392), .Z(N144) );
  GTECH_XOR2 U379 ( .A(n394), .B(n395), .Z(n392) );
  GTECH_OA21 U380 ( .A(n380), .B(n381), .C(n382), .Z(n395) );
  GTECH_OAI21 U381 ( .A(n396), .B(n397), .C(n398), .Z(n382) );
  GTECH_XOR4 U382 ( .A(n378), .B(n387), .C(n388), .D(n376), .Z(n394) );
  GTECH_XNOR3 U383 ( .A(n399), .B(n400), .C(n401), .Z(n376) );
  GTECH_NOT U384 ( .A(n385), .Z(n401) );
  GTECH_NAND3 U385 ( .A(I_b[2]), .B(I_a[1]), .C(n402), .Z(n385) );
  GTECH_NOT U386 ( .A(n384), .Z(n400) );
  GTECH_OR_NOT U387 ( .A(n276), .B(I_b[3]), .Z(n384) );
  GTECH_NOT U388 ( .A(n383), .Z(n399) );
  GTECH_OR_NOT U389 ( .A(n238), .B(I_b[2]), .Z(n383) );
  GTECH_OR_NOT U390 ( .A(n341), .B(I_a[4]), .Z(n388) );
  GTECH_NOT U391 ( .A(I_b[0]), .Z(n341) );
  GTECH_NOT U392 ( .A(n379), .Z(n387) );
  GTECH_OAI21 U393 ( .A(n403), .B(n404), .C(n405), .Z(n379) );
  GTECH_OAI21 U394 ( .A(n406), .B(n407), .C(n408), .Z(n405) );
  GTECH_NOT U395 ( .A(n409), .Z(n378) );
  GTECH_OR_NOT U396 ( .A(n340), .B(I_a[3]), .Z(n409) );
  GTECH_AND2 U397 ( .A(I_b[4]), .B(I_a[0]), .Z(n393) );
  GTECH_XNOR3 U398 ( .A(n398), .B(n381), .C(n397), .Z(N143) );
  GTECH_NOT U399 ( .A(n380), .Z(n397) );
  GTECH_XOR2 U400 ( .A(n410), .B(n402), .Z(n380) );
  GTECH_NOT U401 ( .A(n411), .Z(n402) );
  GTECH_OR_NOT U402 ( .A(n320), .B(I_b[3]), .Z(n411) );
  GTECH_NOT U403 ( .A(I_a[0]), .Z(n320) );
  GTECH_OR_NOT U404 ( .A(n276), .B(I_b[2]), .Z(n410) );
  GTECH_NOT U405 ( .A(I_a[1]), .Z(n276) );
  GTECH_NOT U406 ( .A(n396), .Z(n381) );
  GTECH_XNOR3 U407 ( .A(n406), .B(n408), .C(n403), .Z(n396) );
  GTECH_NOT U408 ( .A(n407), .Z(n403) );
  GTECH_OAI21 U409 ( .A(n412), .B(n413), .C(n414), .Z(n407) );
  GTECH_NOT U410 ( .A(n415), .Z(n408) );
  GTECH_OR_NOT U411 ( .A(n238), .B(I_b[1]), .Z(n415) );
  GTECH_NOT U412 ( .A(n404), .Z(n406) );
  GTECH_OR_NOT U413 ( .A(n201), .B(I_b[0]), .Z(n404) );
  GTECH_NOT U414 ( .A(I_a[3]), .Z(n201) );
  GTECH_NOT U415 ( .A(n416), .Z(n398) );
  GTECH_NAND3 U416 ( .A(I_a[0]), .B(n417), .C(I_b[2]), .Z(n416) );
  GTECH_XOR2 U417 ( .A(n418), .B(n417), .Z(N142) );
  GTECH_NOT U418 ( .A(n419), .Z(n417) );
  GTECH_XNOR3 U419 ( .A(n420), .B(n421), .C(n422), .Z(n419) );
  GTECH_NOT U420 ( .A(n414), .Z(n422) );
  GTECH_NAND3 U421 ( .A(n423), .B(I_b[0]), .C(I_a[1]), .Z(n414) );
  GTECH_NOT U422 ( .A(n412), .Z(n421) );
  GTECH_OR_NOT U423 ( .A(n340), .B(I_a[1]), .Z(n412) );
  GTECH_NOT U424 ( .A(n413), .Z(n420) );
  GTECH_OR_NOT U425 ( .A(n238), .B(I_b[0]), .Z(n413) );
  GTECH_NOT U426 ( .A(I_a[2]), .Z(n238) );
  GTECH_AND2 U427 ( .A(I_b[2]), .B(I_a[0]), .Z(n418) );
  GTECH_XOR2 U428 ( .A(n423), .B(n424), .Z(N141) );
  GTECH_AND2 U429 ( .A(I_a[1]), .B(I_b[0]), .Z(n424) );
  GTECH_NOT U430 ( .A(n425), .Z(n423) );
  GTECH_OR_NOT U431 ( .A(n340), .B(I_a[0]), .Z(n425) );
  GTECH_NOT U432 ( .A(I_b[1]), .Z(n340) );
  GTECH_AND2 U433 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

