
module array_multiplier16 ( clk, I_reset_n, I_valid, I_a, I_b, O_valid, O_c );
  input [7:0] I_a;
  input [7:0] I_b;
  output [15:0] O_c;
  input clk, I_reset_n, I_valid;
  output O_valid;
  wire   N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409;

  GTECH_FD2 O_valid_reg ( .D(I_valid), .CP(clk), .CD(I_reset_n), .Q(O_valid)
         );
  GTECH_FD2 O_c_reg_15_ ( .D(N155), .CP(clk), .CD(I_reset_n), .Q(O_c[15]) );
  GTECH_FD2 O_c_reg_14_ ( .D(N154), .CP(clk), .CD(I_reset_n), .Q(O_c[14]) );
  GTECH_FD2 O_c_reg_13_ ( .D(N153), .CP(clk), .CD(I_reset_n), .Q(O_c[13]) );
  GTECH_FD2 O_c_reg_12_ ( .D(N152), .CP(clk), .CD(I_reset_n), .Q(O_c[12]) );
  GTECH_FD2 O_c_reg_11_ ( .D(N151), .CP(clk), .CD(I_reset_n), .Q(O_c[11]) );
  GTECH_FD2 O_c_reg_10_ ( .D(N150), .CP(clk), .CD(I_reset_n), .Q(O_c[10]) );
  GTECH_FD2 O_c_reg_9_ ( .D(N149), .CP(clk), .CD(I_reset_n), .Q(O_c[9]) );
  GTECH_FD2 O_c_reg_8_ ( .D(N148), .CP(clk), .CD(I_reset_n), .Q(O_c[8]) );
  GTECH_FD2 O_c_reg_7_ ( .D(N147), .CP(clk), .CD(I_reset_n), .Q(O_c[7]) );
  GTECH_FD2 O_c_reg_6_ ( .D(N146), .CP(clk), .CD(I_reset_n), .Q(O_c[6]) );
  GTECH_FD2 O_c_reg_5_ ( .D(N145), .CP(clk), .CD(I_reset_n), .Q(O_c[5]) );
  GTECH_FD2 O_c_reg_4_ ( .D(N144), .CP(clk), .CD(I_reset_n), .Q(O_c[4]) );
  GTECH_FD2 O_c_reg_3_ ( .D(N143), .CP(clk), .CD(I_reset_n), .Q(O_c[3]) );
  GTECH_FD2 O_c_reg_2_ ( .D(N142), .CP(clk), .CD(I_reset_n), .Q(O_c[2]) );
  GTECH_FD2 O_c_reg_1_ ( .D(N141), .CP(clk), .CD(I_reset_n), .Q(O_c[1]) );
  GTECH_FD2 O_c_reg_0_ ( .D(N140), .CP(clk), .CD(I_reset_n), .Q(O_c[0]) );
  GTECH_NOT U75 ( .A(n83), .Z(N155) );
  GTECH_AOI222 U76 ( .A(n84), .B(n85), .C(n86), .D(n87), .E(n88), .F(n89), .Z(
        n83) );
  GTECH_NOT U77 ( .A(n90), .Z(n88) );
  GTECH_XOR2 U78 ( .A(n84), .B(n85), .Z(N154) );
  GTECH_NOT U79 ( .A(n91), .Z(n85) );
  GTECH_XOR2 U80 ( .A(n86), .B(n92), .Z(n91) );
  GTECH_NOT U81 ( .A(n87), .Z(n92) );
  GTECH_OAI22 U82 ( .A(n93), .B(n94), .C(n95), .D(n96), .Z(n87) );
  GTECH_AND2 U83 ( .A(n93), .B(n94), .Z(n95) );
  GTECH_XOR2 U84 ( .A(n90), .B(n97), .Z(n86) );
  GTECH_NOT U85 ( .A(n89), .Z(n97) );
  GTECH_OAI22 U86 ( .A(n98), .B(n99), .C(n100), .D(n101), .Z(n89) );
  GTECH_AND2 U87 ( .A(n98), .B(n99), .Z(n100) );
  GTECH_NAND2 U88 ( .A(I_b[7]), .B(I_a[7]), .Z(n90) );
  GTECH_NOT U89 ( .A(n102), .Z(n84) );
  GTECH_NAND2 U90 ( .A(n103), .B(n104), .Z(n102) );
  GTECH_XOR2 U91 ( .A(n104), .B(n103), .Z(N153) );
  GTECH_NOT U92 ( .A(n105), .Z(n103) );
  GTECH_XNOR3 U93 ( .A(n106), .B(n93), .C(n96), .Z(n105) );
  GTECH_NOT U94 ( .A(n107), .Z(n96) );
  GTECH_XNOR3 U95 ( .A(n108), .B(n109), .C(n98), .Z(n107) );
  GTECH_OA21 U96 ( .A(n110), .B(n111), .C(n112), .Z(n98) );
  GTECH_AO21 U97 ( .A(n110), .B(n111), .C(n113), .Z(n112) );
  GTECH_NOT U98 ( .A(n101), .Z(n109) );
  GTECH_NAND2 U99 ( .A(I_b[7]), .B(I_a[6]), .Z(n101) );
  GTECH_NOT U100 ( .A(n99), .Z(n108) );
  GTECH_NAND2 U101 ( .A(I_a[7]), .B(I_b[6]), .Z(n99) );
  GTECH_ADD_ABC U102 ( .A(n114), .B(n115), .C(n116), .COUT(n93) );
  GTECH_NOT U103 ( .A(n117), .Z(n116) );
  GTECH_XOR2 U104 ( .A(n118), .B(n119), .Z(n115) );
  GTECH_AND2 U105 ( .A(I_a[7]), .B(I_b[5]), .Z(n119) );
  GTECH_NOT U106 ( .A(n94), .Z(n106) );
  GTECH_NAND2 U107 ( .A(I_a[7]), .B(n120), .Z(n94) );
  GTECH_NOT U108 ( .A(n121), .Z(n104) );
  GTECH_NAND2 U109 ( .A(n122), .B(n123), .Z(n121) );
  GTECH_NOT U110 ( .A(n124), .Z(n123) );
  GTECH_XOR2 U111 ( .A(n124), .B(n125), .Z(N152) );
  GTECH_NOT U112 ( .A(n122), .Z(n125) );
  GTECH_XOR4 U113 ( .A(n126), .B(n118), .C(n117), .D(n114), .Z(n122) );
  GTECH_ADD_ABC U114 ( .A(n127), .B(n128), .C(n129), .COUT(n114) );
  GTECH_XNOR3 U115 ( .A(n130), .B(n131), .C(n132), .Z(n128) );
  GTECH_XNOR3 U116 ( .A(n133), .B(n134), .C(n110), .Z(n117) );
  GTECH_OA21 U117 ( .A(n135), .B(n136), .C(n137), .Z(n110) );
  GTECH_AO21 U118 ( .A(n135), .B(n136), .C(n138), .Z(n137) );
  GTECH_NOT U119 ( .A(n113), .Z(n134) );
  GTECH_NAND2 U120 ( .A(I_b[7]), .B(I_a[5]), .Z(n113) );
  GTECH_NOT U121 ( .A(n111), .Z(n133) );
  GTECH_NAND2 U122 ( .A(I_b[6]), .B(I_a[6]), .Z(n111) );
  GTECH_NOT U123 ( .A(n120), .Z(n118) );
  GTECH_OAI22 U124 ( .A(n139), .B(n140), .C(n141), .D(n142), .Z(n120) );
  GTECH_AND2 U125 ( .A(n139), .B(n140), .Z(n141) );
  GTECH_AND2 U126 ( .A(I_a[7]), .B(I_b[5]), .Z(n126) );
  GTECH_ADD_ABC U127 ( .A(n143), .B(n144), .C(n145), .COUT(n124) );
  GTECH_OA22 U128 ( .A(n146), .B(n147), .C(n148), .D(n149), .Z(n144) );
  GTECH_OA21 U129 ( .A(n150), .B(n151), .C(n152), .Z(n143) );
  GTECH_AO21 U130 ( .A(n150), .B(n151), .C(n153), .Z(n152) );
  GTECH_XNOR3 U131 ( .A(n154), .B(n145), .C(n155), .Z(N151) );
  GTECH_OA21 U132 ( .A(n150), .B(n151), .C(n156), .Z(n155) );
  GTECH_AO21 U133 ( .A(n150), .B(n151), .C(n153), .Z(n156) );
  GTECH_NOT U134 ( .A(n157), .Z(n153) );
  GTECH_XOR2 U135 ( .A(n127), .B(n158), .Z(n145) );
  GTECH_XOR4 U136 ( .A(n131), .B(n139), .C(n129), .D(n130), .Z(n158) );
  GTECH_NOT U137 ( .A(n140), .Z(n130) );
  GTECH_NAND2 U138 ( .A(I_a[7]), .B(I_b[4]), .Z(n140) );
  GTECH_NOT U139 ( .A(n159), .Z(n129) );
  GTECH_XNOR3 U140 ( .A(n160), .B(n161), .C(n135), .Z(n159) );
  GTECH_OA21 U141 ( .A(n162), .B(n163), .C(n164), .Z(n135) );
  GTECH_AO21 U142 ( .A(n162), .B(n163), .C(n165), .Z(n164) );
  GTECH_NOT U143 ( .A(n138), .Z(n161) );
  GTECH_NAND2 U144 ( .A(I_b[7]), .B(I_a[4]), .Z(n138) );
  GTECH_NOT U145 ( .A(n136), .Z(n160) );
  GTECH_NAND2 U146 ( .A(I_b[6]), .B(I_a[5]), .Z(n136) );
  GTECH_NOT U147 ( .A(n132), .Z(n139) );
  GTECH_OAI22 U148 ( .A(n166), .B(n167), .C(n168), .D(n169), .Z(n132) );
  GTECH_AND2 U149 ( .A(n166), .B(n167), .Z(n168) );
  GTECH_NOT U150 ( .A(n142), .Z(n131) );
  GTECH_NAND2 U151 ( .A(I_a[6]), .B(I_b[5]), .Z(n142) );
  GTECH_ADD_ABC U152 ( .A(n170), .B(n171), .C(n172), .COUT(n127) );
  GTECH_NOT U153 ( .A(n173), .Z(n172) );
  GTECH_XNOR3 U154 ( .A(n174), .B(n175), .C(n176), .Z(n171) );
  GTECH_OA22 U155 ( .A(n146), .B(n147), .C(n148), .D(n149), .Z(n154) );
  GTECH_NOT U156 ( .A(n177), .Z(n149) );
  GTECH_NOT U157 ( .A(I_a[7]), .Z(n147) );
  GTECH_XNOR3 U158 ( .A(n150), .B(n178), .C(n157), .Z(N150) );
  GTECH_XOR2 U159 ( .A(n179), .B(n170), .Z(n157) );
  GTECH_ADD_ABC U160 ( .A(n180), .B(n181), .C(n182), .COUT(n170) );
  GTECH_NOT U161 ( .A(n183), .Z(n182) );
  GTECH_XNOR3 U162 ( .A(n184), .B(n185), .C(n186), .Z(n181) );
  GTECH_XOR4 U163 ( .A(n175), .B(n166), .C(n173), .D(n174), .Z(n179) );
  GTECH_NOT U164 ( .A(n167), .Z(n174) );
  GTECH_NAND2 U165 ( .A(I_a[6]), .B(I_b[4]), .Z(n167) );
  GTECH_XNOR3 U166 ( .A(n187), .B(n188), .C(n162), .Z(n173) );
  GTECH_OA21 U167 ( .A(n189), .B(n190), .C(n191), .Z(n162) );
  GTECH_AO21 U168 ( .A(n189), .B(n190), .C(n192), .Z(n191) );
  GTECH_NOT U169 ( .A(n165), .Z(n188) );
  GTECH_NAND2 U170 ( .A(I_b[7]), .B(I_a[3]), .Z(n165) );
  GTECH_NOT U171 ( .A(n163), .Z(n187) );
  GTECH_NAND2 U172 ( .A(I_b[6]), .B(I_a[4]), .Z(n163) );
  GTECH_NOT U173 ( .A(n176), .Z(n166) );
  GTECH_OAI22 U174 ( .A(n193), .B(n194), .C(n195), .D(n196), .Z(n176) );
  GTECH_AND2 U175 ( .A(n193), .B(n194), .Z(n195) );
  GTECH_NOT U176 ( .A(n169), .Z(n175) );
  GTECH_NAND2 U177 ( .A(I_a[5]), .B(I_b[5]), .Z(n169) );
  GTECH_NOT U178 ( .A(n151), .Z(n178) );
  GTECH_XOR2 U179 ( .A(n177), .B(n148), .Z(n151) );
  GTECH_OA21 U180 ( .A(n197), .B(n198), .C(n199), .Z(n148) );
  GTECH_AO21 U181 ( .A(n197), .B(n198), .C(n200), .Z(n199) );
  GTECH_XOR2 U182 ( .A(n201), .B(n146), .Z(n177) );
  GTECH_OA21 U183 ( .A(n202), .B(n203), .C(n204), .Z(n146) );
  GTECH_AO21 U184 ( .A(n202), .B(n203), .C(n205), .Z(n204) );
  GTECH_NAND2 U185 ( .A(I_a[7]), .B(I_b[3]), .Z(n201) );
  GTECH_AOI2N2 U186 ( .A(n206), .B(n207), .C(n208), .D(n209), .Z(n150) );
  GTECH_NAND2 U187 ( .A(n208), .B(n209), .Z(n207) );
  GTECH_XNOR3 U188 ( .A(n208), .B(n210), .C(n206), .Z(N149) );
  GTECH_XOR2 U189 ( .A(n211), .B(n180), .Z(n206) );
  GTECH_ADD_ABC U190 ( .A(n212), .B(n213), .C(n214), .COUT(n180) );
  GTECH_XNOR3 U191 ( .A(n215), .B(n216), .C(n217), .Z(n213) );
  GTECH_OA21 U192 ( .A(n218), .B(n219), .C(n220), .Z(n212) );
  GTECH_AO21 U193 ( .A(n218), .B(n219), .C(n221), .Z(n220) );
  GTECH_XOR4 U194 ( .A(n185), .B(n193), .C(n183), .D(n184), .Z(n211) );
  GTECH_NOT U195 ( .A(n194), .Z(n184) );
  GTECH_NAND2 U196 ( .A(I_a[5]), .B(I_b[4]), .Z(n194) );
  GTECH_XNOR3 U197 ( .A(n222), .B(n223), .C(n189), .Z(n183) );
  GTECH_NOT U198 ( .A(n224), .Z(n189) );
  GTECH_AO21 U199 ( .A(n225), .B(n226), .C(n227), .Z(n224) );
  GTECH_NOT U200 ( .A(n192), .Z(n223) );
  GTECH_NAND2 U201 ( .A(I_b[7]), .B(I_a[2]), .Z(n192) );
  GTECH_NOT U202 ( .A(n190), .Z(n222) );
  GTECH_NAND2 U203 ( .A(I_b[6]), .B(I_a[3]), .Z(n190) );
  GTECH_NOT U204 ( .A(n186), .Z(n193) );
  GTECH_OAI22 U205 ( .A(n228), .B(n229), .C(n230), .D(n231), .Z(n186) );
  GTECH_AND2 U206 ( .A(n228), .B(n229), .Z(n230) );
  GTECH_NOT U207 ( .A(n196), .Z(n185) );
  GTECH_NAND2 U208 ( .A(I_b[5]), .B(I_a[4]), .Z(n196) );
  GTECH_NOT U209 ( .A(n209), .Z(n210) );
  GTECH_XNOR3 U210 ( .A(n232), .B(n197), .C(n200), .Z(n209) );
  GTECH_NOT U211 ( .A(n233), .Z(n200) );
  GTECH_XNOR3 U212 ( .A(n234), .B(n235), .C(n202), .Z(n233) );
  GTECH_OA21 U213 ( .A(n236), .B(n237), .C(n238), .Z(n202) );
  GTECH_AO21 U214 ( .A(n236), .B(n237), .C(n239), .Z(n238) );
  GTECH_NOT U215 ( .A(n205), .Z(n235) );
  GTECH_NAND2 U216 ( .A(I_a[6]), .B(I_b[3]), .Z(n205) );
  GTECH_NOT U217 ( .A(n203), .Z(n234) );
  GTECH_NAND2 U218 ( .A(I_a[7]), .B(I_b[2]), .Z(n203) );
  GTECH_ADD_ABC U219 ( .A(n240), .B(n241), .C(n242), .COUT(n197) );
  GTECH_NOT U220 ( .A(n243), .Z(n242) );
  GTECH_XOR2 U221 ( .A(n244), .B(n245), .Z(n241) );
  GTECH_AND2 U222 ( .A(I_a[7]), .B(I_b[1]), .Z(n245) );
  GTECH_NOT U223 ( .A(n198), .Z(n232) );
  GTECH_NAND2 U224 ( .A(I_a[7]), .B(n246), .Z(n198) );
  GTECH_ADD_ABC U225 ( .A(n247), .B(n248), .C(n249), .COUT(n208) );
  GTECH_XNOR3 U226 ( .A(n240), .B(n250), .C(n243), .Z(n248) );
  GTECH_XOR2 U227 ( .A(n251), .B(n247), .Z(N148) );
  GTECH_ADD_ABC U228 ( .A(n252), .B(n253), .C(n254), .COUT(n247) );
  GTECH_NOT U229 ( .A(n255), .Z(n254) );
  GTECH_XNOR3 U230 ( .A(n256), .B(n257), .C(n258), .Z(n253) );
  GTECH_XOR4 U231 ( .A(n250), .B(n240), .C(n243), .D(n249), .Z(n251) );
  GTECH_XOR2 U232 ( .A(n259), .B(n260), .Z(n249) );
  GTECH_XOR4 U233 ( .A(n216), .B(n228), .C(n214), .D(n215), .Z(n260) );
  GTECH_NOT U234 ( .A(n229), .Z(n215) );
  GTECH_NAND2 U235 ( .A(I_b[4]), .B(I_a[4]), .Z(n229) );
  GTECH_XNOR3 U236 ( .A(n226), .B(n225), .C(n227), .Z(n214) );
  GTECH_NOT U237 ( .A(n261), .Z(n227) );
  GTECH_NAND3 U238 ( .A(I_b[6]), .B(I_a[1]), .C(n262), .Z(n261) );
  GTECH_NOT U239 ( .A(n263), .Z(n225) );
  GTECH_NAND2 U240 ( .A(I_b[7]), .B(I_a[1]), .Z(n263) );
  GTECH_NOT U241 ( .A(n264), .Z(n226) );
  GTECH_NAND2 U242 ( .A(I_b[6]), .B(I_a[2]), .Z(n264) );
  GTECH_NOT U243 ( .A(n217), .Z(n228) );
  GTECH_OAI22 U244 ( .A(n265), .B(n266), .C(n267), .D(n268), .Z(n217) );
  GTECH_AND2 U245 ( .A(n265), .B(n266), .Z(n267) );
  GTECH_NOT U246 ( .A(n231), .Z(n216) );
  GTECH_NAND2 U247 ( .A(I_b[5]), .B(I_a[3]), .Z(n231) );
  GTECH_OA21 U248 ( .A(n218), .B(n219), .C(n269), .Z(n259) );
  GTECH_AO21 U249 ( .A(n218), .B(n219), .C(n221), .Z(n269) );
  GTECH_XNOR3 U250 ( .A(n270), .B(n271), .C(n236), .Z(n243) );
  GTECH_OA21 U251 ( .A(n272), .B(n273), .C(n274), .Z(n236) );
  GTECH_AO21 U252 ( .A(n272), .B(n273), .C(n275), .Z(n274) );
  GTECH_NOT U253 ( .A(n239), .Z(n271) );
  GTECH_NAND2 U254 ( .A(I_a[5]), .B(I_b[3]), .Z(n239) );
  GTECH_NOT U255 ( .A(n237), .Z(n270) );
  GTECH_NAND2 U256 ( .A(I_a[6]), .B(I_b[2]), .Z(n237) );
  GTECH_ADD_ABC U257 ( .A(n256), .B(n276), .C(n277), .COUT(n240) );
  GTECH_XNOR3 U258 ( .A(n278), .B(n279), .C(n280), .Z(n276) );
  GTECH_XOR2 U259 ( .A(n281), .B(n244), .Z(n250) );
  GTECH_NOT U260 ( .A(n246), .Z(n244) );
  GTECH_OAI22 U261 ( .A(n282), .B(n283), .C(n284), .D(n285), .Z(n246) );
  GTECH_AND2 U262 ( .A(n282), .B(n283), .Z(n284) );
  GTECH_AND2 U263 ( .A(I_a[7]), .B(I_b[1]), .Z(n281) );
  GTECH_XOR2 U264 ( .A(n286), .B(n252), .Z(N147) );
  GTECH_ADD_ABC U265 ( .A(n287), .B(n288), .C(n289), .COUT(n252) );
  GTECH_XNOR3 U266 ( .A(n290), .B(n291), .C(n292), .Z(n288) );
  GTECH_OA21 U267 ( .A(n293), .B(n294), .C(n295), .Z(n287) );
  GTECH_AO21 U268 ( .A(n293), .B(n294), .C(n296), .Z(n295) );
  GTECH_XOR4 U269 ( .A(n257), .B(n277), .C(n255), .D(n256), .Z(n286) );
  GTECH_ADD_ABC U270 ( .A(n290), .B(n297), .C(n298), .COUT(n256) );
  GTECH_NOT U271 ( .A(n292), .Z(n298) );
  GTECH_XNOR3 U272 ( .A(n299), .B(n300), .C(n301), .Z(n297) );
  GTECH_XNOR3 U273 ( .A(n302), .B(n219), .C(n303), .Z(n255) );
  GTECH_NOT U274 ( .A(n218), .Z(n303) );
  GTECH_XOR2 U275 ( .A(n304), .B(n262), .Z(n218) );
  GTECH_NOT U276 ( .A(n305), .Z(n262) );
  GTECH_NAND2 U277 ( .A(I_b[7]), .B(I_a[0]), .Z(n305) );
  GTECH_NAND2 U278 ( .A(I_b[6]), .B(I_a[1]), .Z(n304) );
  GTECH_NOT U279 ( .A(n306), .Z(n219) );
  GTECH_XNOR3 U280 ( .A(n307), .B(n308), .C(n265), .Z(n306) );
  GTECH_NOT U281 ( .A(n309), .Z(n265) );
  GTECH_AO21 U282 ( .A(n310), .B(n311), .C(n312), .Z(n309) );
  GTECH_NOT U283 ( .A(n268), .Z(n308) );
  GTECH_NAND2 U284 ( .A(I_b[5]), .B(I_a[2]), .Z(n268) );
  GTECH_NOT U285 ( .A(n266), .Z(n307) );
  GTECH_NAND2 U286 ( .A(I_b[4]), .B(I_a[3]), .Z(n266) );
  GTECH_NOT U287 ( .A(n221), .Z(n302) );
  GTECH_NAND3 U288 ( .A(I_a[0]), .B(n313), .C(I_b[6]), .Z(n221) );
  GTECH_NOT U289 ( .A(n314), .Z(n313) );
  GTECH_NOT U290 ( .A(n258), .Z(n277) );
  GTECH_XNOR3 U291 ( .A(n315), .B(n316), .C(n272), .Z(n258) );
  GTECH_OA21 U292 ( .A(n317), .B(n318), .C(n319), .Z(n272) );
  GTECH_AO21 U293 ( .A(n317), .B(n318), .C(n320), .Z(n319) );
  GTECH_NOT U294 ( .A(n275), .Z(n316) );
  GTECH_NAND2 U295 ( .A(I_b[3]), .B(I_a[4]), .Z(n275) );
  GTECH_NOT U296 ( .A(n273), .Z(n315) );
  GTECH_NAND2 U297 ( .A(I_a[5]), .B(I_b[2]), .Z(n273) );
  GTECH_NOT U298 ( .A(n321), .Z(n257) );
  GTECH_XNOR3 U299 ( .A(n278), .B(n279), .C(n282), .Z(n321) );
  GTECH_NOT U300 ( .A(n280), .Z(n282) );
  GTECH_OAI22 U301 ( .A(n322), .B(n323), .C(n324), .D(n325), .Z(n280) );
  GTECH_AND2 U302 ( .A(n322), .B(n323), .Z(n324) );
  GTECH_NOT U303 ( .A(n285), .Z(n279) );
  GTECH_NAND2 U304 ( .A(I_a[6]), .B(I_b[1]), .Z(n285) );
  GTECH_NOT U305 ( .A(n283), .Z(n278) );
  GTECH_NAND2 U306 ( .A(I_a[7]), .B(I_b[0]), .Z(n283) );
  GTECH_XOR2 U307 ( .A(n326), .B(n327), .Z(N146) );
  GTECH_OA21 U308 ( .A(n293), .B(n294), .C(n328), .Z(n327) );
  GTECH_AO21 U309 ( .A(n293), .B(n294), .C(n296), .Z(n328) );
  GTECH_XOR4 U310 ( .A(n291), .B(n290), .C(n292), .D(n289), .Z(n326) );
  GTECH_XOR2 U311 ( .A(n314), .B(n329), .Z(n289) );
  GTECH_AND2 U312 ( .A(I_b[6]), .B(I_a[0]), .Z(n329) );
  GTECH_XNOR3 U313 ( .A(n311), .B(n310), .C(n312), .Z(n314) );
  GTECH_NOT U314 ( .A(n330), .Z(n312) );
  GTECH_NAND3 U315 ( .A(I_b[4]), .B(I_a[1]), .C(n331), .Z(n330) );
  GTECH_NOT U316 ( .A(n332), .Z(n310) );
  GTECH_NAND2 U317 ( .A(I_b[5]), .B(I_a[1]), .Z(n332) );
  GTECH_NOT U318 ( .A(n333), .Z(n311) );
  GTECH_NAND2 U319 ( .A(I_b[4]), .B(I_a[2]), .Z(n333) );
  GTECH_XNOR3 U320 ( .A(n334), .B(n335), .C(n317), .Z(n292) );
  GTECH_OA21 U321 ( .A(n336), .B(n337), .C(n338), .Z(n317) );
  GTECH_AO21 U322 ( .A(n336), .B(n337), .C(n339), .Z(n338) );
  GTECH_NOT U323 ( .A(n320), .Z(n335) );
  GTECH_NAND2 U324 ( .A(I_b[3]), .B(I_a[3]), .Z(n320) );
  GTECH_NOT U325 ( .A(n318), .Z(n334) );
  GTECH_NAND2 U326 ( .A(I_b[2]), .B(I_a[4]), .Z(n318) );
  GTECH_ADD_ABC U327 ( .A(n340), .B(n341), .C(n342), .COUT(n290) );
  GTECH_XNOR3 U328 ( .A(n343), .B(n344), .C(n345), .Z(n341) );
  GTECH_NOT U329 ( .A(n346), .Z(n291) );
  GTECH_XNOR3 U330 ( .A(n299), .B(n300), .C(n322), .Z(n346) );
  GTECH_NOT U331 ( .A(n301), .Z(n322) );
  GTECH_OAI22 U332 ( .A(n347), .B(n348), .C(n349), .D(n350), .Z(n301) );
  GTECH_AND2 U333 ( .A(n347), .B(n348), .Z(n349) );
  GTECH_NOT U334 ( .A(n325), .Z(n300) );
  GTECH_NAND2 U335 ( .A(I_a[5]), .B(I_b[1]), .Z(n325) );
  GTECH_NOT U336 ( .A(n323), .Z(n299) );
  GTECH_NAND2 U337 ( .A(I_a[6]), .B(I_b[0]), .Z(n323) );
  GTECH_XNOR3 U338 ( .A(n351), .B(n294), .C(n352), .Z(N145) );
  GTECH_NOT U339 ( .A(n293), .Z(n352) );
  GTECH_XOR2 U340 ( .A(n353), .B(n331), .Z(n293) );
  GTECH_NOT U341 ( .A(n354), .Z(n331) );
  GTECH_NAND2 U342 ( .A(I_b[5]), .B(I_a[0]), .Z(n354) );
  GTECH_NAND2 U343 ( .A(I_b[4]), .B(I_a[1]), .Z(n353) );
  GTECH_XOR2 U344 ( .A(n340), .B(n355), .Z(n294) );
  GTECH_XOR4 U345 ( .A(n344), .B(n347), .C(n342), .D(n343), .Z(n355) );
  GTECH_NOT U346 ( .A(n348), .Z(n343) );
  GTECH_NAND2 U347 ( .A(I_a[5]), .B(I_b[0]), .Z(n348) );
  GTECH_NOT U348 ( .A(n356), .Z(n342) );
  GTECH_XNOR3 U349 ( .A(n357), .B(n358), .C(n336), .Z(n356) );
  GTECH_NOT U350 ( .A(n359), .Z(n336) );
  GTECH_AO21 U351 ( .A(n360), .B(n361), .C(n362), .Z(n359) );
  GTECH_NOT U352 ( .A(n339), .Z(n358) );
  GTECH_NAND2 U353 ( .A(I_b[3]), .B(I_a[2]), .Z(n339) );
  GTECH_NOT U354 ( .A(n337), .Z(n357) );
  GTECH_NAND2 U355 ( .A(I_b[2]), .B(I_a[3]), .Z(n337) );
  GTECH_NOT U356 ( .A(n345), .Z(n347) );
  GTECH_OAI22 U357 ( .A(n363), .B(n364), .C(n365), .D(n366), .Z(n345) );
  GTECH_AND2 U358 ( .A(n363), .B(n364), .Z(n365) );
  GTECH_NOT U359 ( .A(n350), .Z(n344) );
  GTECH_NAND2 U360 ( .A(I_a[4]), .B(I_b[1]), .Z(n350) );
  GTECH_ADD_ABC U361 ( .A(n367), .B(n368), .C(n369), .COUT(n340) );
  GTECH_XNOR3 U362 ( .A(n370), .B(n371), .C(n372), .Z(n368) );
  GTECH_NOT U363 ( .A(n364), .Z(n370) );
  GTECH_OA21 U364 ( .A(n373), .B(n374), .C(n375), .Z(n367) );
  GTECH_AO21 U365 ( .A(n373), .B(n374), .C(n376), .Z(n375) );
  GTECH_NOT U366 ( .A(n296), .Z(n351) );
  GTECH_NAND3 U367 ( .A(I_a[0]), .B(n377), .C(I_b[4]), .Z(n296) );
  GTECH_XOR2 U368 ( .A(n378), .B(n377), .Z(N144) );
  GTECH_XOR2 U369 ( .A(n379), .B(n380), .Z(n377) );
  GTECH_OA21 U370 ( .A(n373), .B(n374), .C(n381), .Z(n380) );
  GTECH_AO21 U371 ( .A(n373), .B(n374), .C(n376), .Z(n381) );
  GTECH_XOR4 U372 ( .A(n371), .B(n363), .C(n364), .D(n369), .Z(n379) );
  GTECH_XNOR3 U373 ( .A(n361), .B(n360), .C(n362), .Z(n369) );
  GTECH_NOT U374 ( .A(n382), .Z(n362) );
  GTECH_NAND3 U375 ( .A(I_b[2]), .B(I_a[1]), .C(n383), .Z(n382) );
  GTECH_NOT U376 ( .A(n384), .Z(n360) );
  GTECH_NAND2 U377 ( .A(I_b[3]), .B(I_a[1]), .Z(n384) );
  GTECH_NOT U378 ( .A(n385), .Z(n361) );
  GTECH_NAND2 U379 ( .A(I_b[2]), .B(I_a[2]), .Z(n385) );
  GTECH_NAND2 U380 ( .A(I_a[4]), .B(I_b[0]), .Z(n364) );
  GTECH_NOT U381 ( .A(n372), .Z(n363) );
  GTECH_OAI22 U382 ( .A(n386), .B(n387), .C(n388), .D(n389), .Z(n372) );
  GTECH_AND2 U383 ( .A(n386), .B(n387), .Z(n388) );
  GTECH_NOT U384 ( .A(n366), .Z(n371) );
  GTECH_NAND2 U385 ( .A(I_a[3]), .B(I_b[1]), .Z(n366) );
  GTECH_AND2 U386 ( .A(I_b[4]), .B(I_a[0]), .Z(n378) );
  GTECH_XNOR3 U387 ( .A(n390), .B(n374), .C(n391), .Z(N143) );
  GTECH_NOT U388 ( .A(n373), .Z(n391) );
  GTECH_XOR2 U389 ( .A(n392), .B(n383), .Z(n373) );
  GTECH_NOT U390 ( .A(n393), .Z(n383) );
  GTECH_NAND2 U391 ( .A(I_b[3]), .B(I_a[0]), .Z(n393) );
  GTECH_NAND2 U392 ( .A(I_b[2]), .B(I_a[1]), .Z(n392) );
  GTECH_NOT U393 ( .A(n394), .Z(n374) );
  GTECH_XNOR3 U394 ( .A(n395), .B(n396), .C(n386), .Z(n394) );
  GTECH_NOT U395 ( .A(n397), .Z(n386) );
  GTECH_AO21 U396 ( .A(n398), .B(n399), .C(n400), .Z(n397) );
  GTECH_NOT U397 ( .A(n389), .Z(n396) );
  GTECH_NAND2 U398 ( .A(I_b[1]), .B(I_a[2]), .Z(n389) );
  GTECH_NOT U399 ( .A(n387), .Z(n395) );
  GTECH_NAND2 U400 ( .A(I_b[0]), .B(I_a[3]), .Z(n387) );
  GTECH_NOT U401 ( .A(n376), .Z(n390) );
  GTECH_NAND3 U402 ( .A(I_a[0]), .B(n401), .C(I_b[2]), .Z(n376) );
  GTECH_XOR2 U403 ( .A(n402), .B(n401), .Z(N142) );
  GTECH_NOT U404 ( .A(n403), .Z(n401) );
  GTECH_XNOR3 U405 ( .A(n398), .B(n399), .C(n400), .Z(n403) );
  GTECH_NOT U406 ( .A(n404), .Z(n400) );
  GTECH_NAND3 U407 ( .A(n405), .B(I_b[0]), .C(I_a[1]), .Z(n404) );
  GTECH_NOT U408 ( .A(n406), .Z(n399) );
  GTECH_NAND2 U409 ( .A(I_a[1]), .B(I_b[1]), .Z(n406) );
  GTECH_NOT U410 ( .A(n407), .Z(n398) );
  GTECH_NAND2 U411 ( .A(I_b[0]), .B(I_a[2]), .Z(n407) );
  GTECH_AND2 U412 ( .A(I_b[2]), .B(I_a[0]), .Z(n402) );
  GTECH_XOR2 U413 ( .A(n405), .B(n408), .Z(N141) );
  GTECH_AND2 U414 ( .A(I_a[1]), .B(I_b[0]), .Z(n408) );
  GTECH_NOT U415 ( .A(n409), .Z(n405) );
  GTECH_NAND2 U416 ( .A(I_a[0]), .B(I_b[1]), .Z(n409) );
  GTECH_AND2 U417 ( .A(I_a[0]), .B(I_b[0]), .Z(N140) );
endmodule

