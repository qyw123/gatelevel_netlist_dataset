
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136;

  GTECH_XOR2 U89 ( .A(n70), .B(n71), .Z(sum[9]) );
  GTECH_XOR2 U90 ( .A(n72), .B(n73), .Z(sum[8]) );
  GTECH_XNOR2 U91 ( .A(n74), .B(n75), .Z(sum[7]) );
  GTECH_OA21 U92 ( .A(n76), .B(n77), .C(n78), .Z(n75) );
  GTECH_XNOR2 U93 ( .A(n76), .B(n79), .Z(sum[6]) );
  GTECH_AOI22 U94 ( .A(n80), .B(n81), .C(b[5]), .D(a[5]), .Z(n76) );
  GTECH_XOR2 U95 ( .A(n81), .B(n80), .Z(sum[5]) );
  GTECH_AO22 U96 ( .A(a[4]), .B(b[4]), .C(n82), .D(n83), .Z(n80) );
  GTECH_XOR2 U97 ( .A(n83), .B(n82), .Z(sum[4]) );
  GTECH_XOR2 U98 ( .A(n84), .B(n85), .Z(sum[3]) );
  GTECH_AO21 U99 ( .A(n86), .B(n87), .C(n88), .Z(n85) );
  GTECH_XOR2 U100 ( .A(n87), .B(n86), .Z(sum[2]) );
  GTECH_AO21 U101 ( .A(n89), .B(n90), .C(n91), .Z(n86) );
  GTECH_XOR2 U102 ( .A(n90), .B(n89), .Z(sum[1]) );
  GTECH_AO22 U103 ( .A(a[0]), .B(b[0]), .C(n92), .D(cin), .Z(n89) );
  GTECH_XOR2 U104 ( .A(n93), .B(n94), .Z(sum[15]) );
  GTECH_AO21 U105 ( .A(n95), .B(n96), .C(n97), .Z(n94) );
  GTECH_XOR2 U106 ( .A(n96), .B(n95), .Z(sum[14]) );
  GTECH_AO21 U107 ( .A(n98), .B(n99), .C(n100), .Z(n95) );
  GTECH_XOR2 U108 ( .A(n99), .B(n98), .Z(sum[13]) );
  GTECH_AO22 U109 ( .A(a[12]), .B(b[12]), .C(cout), .D(n101), .Z(n98) );
  GTECH_XOR2 U110 ( .A(n101), .B(cout), .Z(sum[12]) );
  GTECH_XNOR2 U111 ( .A(n102), .B(n103), .Z(sum[11]) );
  GTECH_OAI21 U112 ( .A(n104), .B(n105), .C(n106), .Z(n102) );
  GTECH_XOR2 U113 ( .A(n105), .B(n104), .Z(sum[10]) );
  GTECH_OA21 U114 ( .A(n71), .B(n70), .C(n107), .Z(n104) );
  GTECH_OA21 U115 ( .A(n73), .B(n72), .C(n108), .Z(n71) );
  GTECH_XOR2 U116 ( .A(cin), .B(n92), .Z(sum[0]) );
  GTECH_OAI21 U117 ( .A(n73), .B(n109), .C(n110), .Z(cout) );
  GTECH_OA21 U118 ( .A(n111), .B(n112), .C(n113), .Z(n73) );
  GTECH_NOT U119 ( .A(n82), .Z(n111) );
  GTECH_OAI21 U120 ( .A(n114), .B(n115), .C(n116), .Z(n82) );
  GTECH_NOT U121 ( .A(cin), .Z(n115) );
  GTECH_NOR3 U122 ( .A(n112), .B(n114), .C(n109), .Z(Pm) );
  GTECH_NAND5 U123 ( .A(n87), .B(n90), .C(n84), .D(n117), .E(n92), .Z(n114) );
  GTECH_XOR2 U124 ( .A(a[0]), .B(b[0]), .Z(n92) );
  GTECH_OAI21 U125 ( .A(n118), .B(n109), .C(n110), .Z(Gm) );
  GTECH_OA21 U126 ( .A(n119), .B(n120), .C(n121), .Z(n110) );
  GTECH_OAI21 U127 ( .A(n97), .B(n122), .C(n93), .Z(n121) );
  GTECH_OA21 U128 ( .A(n100), .B(n123), .C(n96), .Z(n122) );
  GTECH_AND3 U129 ( .A(a[12]), .B(n99), .C(b[12]), .Z(n123) );
  GTECH_AND2 U130 ( .A(b[13]), .B(a[13]), .Z(n100) );
  GTECH_NOT U131 ( .A(a[15]), .Z(n120) );
  GTECH_NAND4 U132 ( .A(n96), .B(n101), .C(n93), .D(n99), .Z(n109) );
  GTECH_XOR2 U133 ( .A(a[13]), .B(b[13]), .Z(n99) );
  GTECH_XNOR2 U134 ( .A(a[15]), .B(n119), .Z(n93) );
  GTECH_NOT U135 ( .A(b[15]), .Z(n119) );
  GTECH_XOR2 U136 ( .A(a[12]), .B(b[12]), .Z(n101) );
  GTECH_OA21 U137 ( .A(b[14]), .B(a[14]), .C(n124), .Z(n96) );
  GTECH_NOT U138 ( .A(n97), .Z(n124) );
  GTECH_AND2 U139 ( .A(b[14]), .B(a[14]), .Z(n97) );
  GTECH_OA21 U140 ( .A(n116), .B(n112), .C(n113), .Z(n118) );
  GTECH_OA21 U141 ( .A(n125), .B(n103), .C(n126), .Z(n113) );
  GTECH_OA21 U142 ( .A(n127), .B(n105), .C(n106), .Z(n125) );
  GTECH_OA21 U143 ( .A(n108), .B(n70), .C(n107), .Z(n127) );
  GTECH_OR4 U144 ( .A(n72), .B(n103), .C(n105), .D(n70), .Z(n112) );
  GTECH_OAI21 U145 ( .A(b[9]), .B(a[9]), .C(n107), .Z(n70) );
  GTECH_NAND2 U146 ( .A(b[9]), .B(a[9]), .Z(n107) );
  GTECH_OAI21 U147 ( .A(b[10]), .B(a[10]), .C(n106), .Z(n105) );
  GTECH_NAND2 U148 ( .A(a[10]), .B(b[10]), .Z(n106) );
  GTECH_OAI21 U149 ( .A(b[11]), .B(a[11]), .C(n126), .Z(n103) );
  GTECH_NAND2 U150 ( .A(b[11]), .B(a[11]), .Z(n126) );
  GTECH_OAI21 U151 ( .A(b[8]), .B(a[8]), .C(n108), .Z(n72) );
  GTECH_NAND2 U152 ( .A(b[8]), .B(a[8]), .Z(n108) );
  GTECH_AOI222 U153 ( .A(a[7]), .B(b[7]), .C(n74), .D(n128), .E(n117), .F(n129), .Z(n116) );
  GTECH_AO21 U154 ( .A(b[3]), .B(a[3]), .C(n130), .Z(n129) );
  GTECH_OA21 U155 ( .A(n131), .B(n88), .C(n84), .Z(n130) );
  GTECH_XOR2 U156 ( .A(a[3]), .B(b[3]), .Z(n84) );
  GTECH_AND2 U157 ( .A(a[2]), .B(b[2]), .Z(n88) );
  GTECH_OA21 U158 ( .A(n132), .B(n91), .C(n87), .Z(n131) );
  GTECH_XOR2 U159 ( .A(a[2]), .B(b[2]), .Z(n87) );
  GTECH_AND2 U160 ( .A(a[1]), .B(b[1]), .Z(n91) );
  GTECH_AND3 U161 ( .A(a[0]), .B(n90), .C(b[0]), .Z(n132) );
  GTECH_XOR2 U162 ( .A(a[1]), .B(b[1]), .Z(n90) );
  GTECH_AND4 U163 ( .A(n79), .B(n83), .C(n74), .D(n81), .Z(n117) );
  GTECH_XOR2 U164 ( .A(a[4]), .B(b[4]), .Z(n83) );
  GTECH_OAI21 U165 ( .A(n133), .B(n77), .C(n78), .Z(n128) );
  GTECH_NOT U166 ( .A(n79), .Z(n77) );
  GTECH_OA21 U167 ( .A(a[6]), .B(b[6]), .C(n78), .Z(n79) );
  GTECH_NAND2 U168 ( .A(b[6]), .B(a[6]), .Z(n78) );
  GTECH_OA21 U169 ( .A(n134), .B(n135), .C(n136), .Z(n133) );
  GTECH_NAND3 U170 ( .A(a[4]), .B(n81), .C(b[4]), .Z(n136) );
  GTECH_XNOR2 U171 ( .A(a[5]), .B(n134), .Z(n81) );
  GTECH_NOT U172 ( .A(a[5]), .Z(n135) );
  GTECH_NOT U173 ( .A(b[5]), .Z(n134) );
  GTECH_XOR2 U174 ( .A(a[7]), .B(b[7]), .Z(n74) );
endmodule

