
module carry_select_adder16 ( a, b, cin, cout, sum );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout;
  wire   n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386;

  GTECH_MUX2 U142 ( .A(n281), .B(n282), .S(n283), .Z(sum[9]) );
  GTECH_XNOR2 U143 ( .A(n284), .B(n285), .Z(n282) );
  GTECH_XNOR2 U144 ( .A(n286), .B(n285), .Z(n281) );
  GTECH_AOI21 U145 ( .A(a[9]), .B(b[9]), .C(n287), .Z(n285) );
  GTECH_NAND2 U146 ( .A(n288), .B(n289), .Z(sum[8]) );
  GTECH_OAI21 U147 ( .A(n290), .B(n284), .C(n283), .Z(n288) );
  GTECH_MUX2 U148 ( .A(n291), .B(n292), .S(n293), .Z(sum[7]) );
  GTECH_XNOR2 U149 ( .A(n294), .B(n295), .Z(n292) );
  GTECH_AND2 U150 ( .A(n296), .B(n297), .Z(n294) );
  GTECH_OAI21 U151 ( .A(b[6]), .B(a[6]), .C(n298), .Z(n297) );
  GTECH_ADD_AB U152 ( .A(n299), .B(n295), .S(n291) );
  GTECH_ADD_AB U153 ( .A(b[7]), .B(a[7]), .S(n295) );
  GTECH_OAI21 U154 ( .A(n300), .B(n296), .C(n301), .Z(sum[6]) );
  GTECH_MUX2 U155 ( .A(n302), .B(n303), .S(b[6]), .Z(n301) );
  GTECH_OR_NOT U156 ( .A(a[6]), .B(n300), .Z(n303) );
  GTECH_ADD_AB U157 ( .A(a[6]), .B(n300), .S(n302) );
  GTECH_AOI21 U158 ( .A(n304), .B(n305), .C(n298), .Z(n300) );
  GTECH_AOI21 U159 ( .A(n306), .B(n307), .C(n308), .Z(n298) );
  GTECH_MUX2 U160 ( .A(n309), .B(n310), .S(n311), .Z(sum[5]) );
  GTECH_AND_NOT U161 ( .A(n306), .B(n308), .Z(n311) );
  GTECH_OAI21 U162 ( .A(a[4]), .B(n305), .C(n312), .Z(n310) );
  GTECH_AO21 U163 ( .A(n305), .B(a[4]), .C(b[4]), .Z(n312) );
  GTECH_OAI21 U164 ( .A(n313), .B(n293), .C(n307), .Z(n309) );
  GTECH_ADD_AB U165 ( .A(n314), .B(n293), .S(sum[4]) );
  GTECH_MUX2 U166 ( .A(n315), .B(n316), .S(cin), .Z(sum[3]) );
  GTECH_ADD_AB U167 ( .A(n317), .B(n318), .S(n316) );
  GTECH_ADD_AB U168 ( .A(n319), .B(n318), .S(n315) );
  GTECH_ADD_AB U169 ( .A(b[3]), .B(a[3]), .S(n318) );
  GTECH_ADD_ABC U170 ( .A(a[2]), .B(n320), .C(b[2]), .COUT(n319) );
  GTECH_MUX2 U171 ( .A(n321), .B(n322), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U172 ( .A(n323), .B(n324), .Z(n322) );
  GTECH_XNOR2 U173 ( .A(n320), .B(n324), .Z(n321) );
  GTECH_XNOR2 U174 ( .A(b[2]), .B(a[2]), .Z(n324) );
  GTECH_OA21 U175 ( .A(n325), .B(n326), .C(n327), .Z(n320) );
  GTECH_MUX2 U176 ( .A(n328), .B(n329), .S(n330), .Z(sum[1]) );
  GTECH_AND_NOT U177 ( .A(n327), .B(n325), .Z(n330) );
  GTECH_OAI21 U178 ( .A(cin), .B(n326), .C(n331), .Z(n329) );
  GTECH_OAI21 U179 ( .A(n332), .B(n333), .C(n334), .Z(n328) );
  GTECH_NOT U180 ( .A(n326), .Z(n334) );
  GTECH_MUX2 U181 ( .A(n335), .B(n336), .S(n337), .Z(sum[15]) );
  GTECH_XNOR2 U182 ( .A(n338), .B(n339), .Z(n336) );
  GTECH_OA21 U183 ( .A(n340), .B(n341), .C(n342), .Z(n338) );
  GTECH_ADD_AB U184 ( .A(n343), .B(n339), .S(n335) );
  GTECH_ADD_AB U185 ( .A(b[15]), .B(a[15]), .S(n339) );
  GTECH_MUX2 U186 ( .A(n344), .B(n345), .S(n346), .Z(sum[14]) );
  GTECH_OA21 U187 ( .A(n347), .B(n337), .C(n341), .Z(n346) );
  GTECH_OA21 U188 ( .A(n348), .B(n349), .C(n350), .Z(n341) );
  GTECH_ADD_AB U189 ( .A(b[14]), .B(a[14]), .S(n345) );
  GTECH_OR_NOT U190 ( .A(n340), .B(n342), .Z(n344) );
  GTECH_MUX2 U191 ( .A(n351), .B(n352), .S(n353), .Z(sum[13]) );
  GTECH_OA21 U192 ( .A(n354), .B(n337), .C(n349), .Z(n353) );
  GTECH_ADD_AB U193 ( .A(b[13]), .B(a[13]), .S(n352) );
  GTECH_OR_NOT U194 ( .A(n348), .B(n350), .Z(n351) );
  GTECH_NAND2 U195 ( .A(n355), .B(n356), .Z(sum[12]) );
  GTECH_OAI21 U196 ( .A(n357), .B(n354), .C(n358), .Z(n355) );
  GTECH_MUX2 U197 ( .A(n359), .B(n360), .S(n283), .Z(sum[11]) );
  GTECH_ADD_AB U198 ( .A(n361), .B(n362), .S(n360) );
  GTECH_XNOR2 U199 ( .A(n363), .B(n362), .Z(n359) );
  GTECH_ADD_AB U200 ( .A(b[11]), .B(a[11]), .S(n362) );
  GTECH_AND2 U201 ( .A(n364), .B(n365), .Z(n363) );
  GTECH_OAI21 U202 ( .A(b[10]), .B(a[10]), .C(n366), .Z(n365) );
  GTECH_OAI21 U203 ( .A(n367), .B(n364), .C(n368), .Z(sum[10]) );
  GTECH_MUX2 U204 ( .A(n369), .B(n370), .S(b[10]), .Z(n368) );
  GTECH_OR_NOT U205 ( .A(a[10]), .B(n367), .Z(n370) );
  GTECH_ADD_AB U206 ( .A(a[10]), .B(n367), .S(n369) );
  GTECH_AOI21 U207 ( .A(n371), .B(n283), .C(n366), .Z(n367) );
  GTECH_OAI2N2 U208 ( .A(n287), .B(n286), .C(a[9]), .D(b[9]), .Z(n366) );
  GTECH_NOT U209 ( .A(n290), .Z(n286) );
  GTECH_XNOR2 U210 ( .A(n333), .B(n372), .Z(sum[0]) );
  GTECH_NOT U211 ( .A(cin), .Z(n333) );
  GTECH_OAI21 U212 ( .A(n337), .B(n373), .C(n356), .Z(cout) );
  GTECH_OR3 U213 ( .A(n357), .B(n354), .C(n358), .Z(n356) );
  GTECH_NOT U214 ( .A(n349), .Z(n357) );
  GTECH_NAND2 U215 ( .A(a[12]), .B(b[12]), .Z(n349) );
  GTECH_AOI21 U216 ( .A(n343), .B(a[15]), .C(n374), .Z(n373) );
  GTECH_OA21 U217 ( .A(a[15]), .B(n343), .C(b[15]), .Z(n374) );
  GTECH_NAND2 U218 ( .A(n375), .B(n342), .Z(n343) );
  GTECH_NAND2 U219 ( .A(a[14]), .B(b[14]), .Z(n342) );
  GTECH_AO21 U220 ( .A(n347), .B(n350), .C(n340), .Z(n375) );
  GTECH_NOR2 U221 ( .A(b[14]), .B(a[14]), .Z(n340) );
  GTECH_NAND2 U222 ( .A(b[13]), .B(a[13]), .Z(n350) );
  GTECH_OR_NOT U223 ( .A(n354), .B(n376), .Z(n347) );
  GTECH_NOT U224 ( .A(n348), .Z(n376) );
  GTECH_NOR2 U225 ( .A(a[13]), .B(b[13]), .Z(n348) );
  GTECH_NOR2 U226 ( .A(b[12]), .B(a[12]), .Z(n354) );
  GTECH_NOT U227 ( .A(n358), .Z(n337) );
  GTECH_OAI21 U228 ( .A(n377), .B(n378), .C(n289), .Z(n358) );
  GTECH_OR3 U229 ( .A(n290), .B(n284), .C(n283), .Z(n289) );
  GTECH_NOT U230 ( .A(n378), .Z(n283) );
  GTECH_AND2 U231 ( .A(b[8]), .B(a[8]), .Z(n290) );
  GTECH_MUX2 U232 ( .A(n379), .B(n314), .S(n293), .Z(n378) );
  GTECH_NOT U233 ( .A(n305), .Z(n293) );
  GTECH_MUX2 U234 ( .A(n372), .B(n380), .S(cin), .Z(n305) );
  GTECH_OA21 U235 ( .A(a[3]), .B(n317), .C(n381), .Z(n380) );
  GTECH_AO21 U236 ( .A(n317), .B(a[3]), .C(b[3]), .Z(n381) );
  GTECH_ADD_ABC U237 ( .A(n323), .B(a[2]), .C(b[2]), .COUT(n317) );
  GTECH_OA21 U238 ( .A(n325), .B(n331), .C(n327), .Z(n323) );
  GTECH_NOT U239 ( .A(n382), .Z(n327) );
  GTECH_NOR2 U240 ( .A(b[1]), .B(a[1]), .Z(n382) );
  GTECH_AND2 U241 ( .A(b[1]), .B(a[1]), .Z(n325) );
  GTECH_AND_NOT U242 ( .A(n331), .B(n326), .Z(n372) );
  GTECH_AND2 U243 ( .A(b[0]), .B(a[0]), .Z(n326) );
  GTECH_NOT U244 ( .A(n332), .Z(n331) );
  GTECH_NOR2 U245 ( .A(b[0]), .B(a[0]), .Z(n332) );
  GTECH_OR_NOT U246 ( .A(n313), .B(n307), .Z(n314) );
  GTECH_NAND2 U247 ( .A(a[4]), .B(b[4]), .Z(n307) );
  GTECH_AOI21 U248 ( .A(n299), .B(a[7]), .C(n383), .Z(n379) );
  GTECH_OA21 U249 ( .A(a[7]), .B(n299), .C(b[7]), .Z(n383) );
  GTECH_NAND2 U250 ( .A(n384), .B(n296), .Z(n299) );
  GTECH_NAND2 U251 ( .A(b[6]), .B(a[6]), .Z(n296) );
  GTECH_OAI21 U252 ( .A(a[6]), .B(b[6]), .C(n304), .Z(n384) );
  GTECH_AOI21 U253 ( .A(n306), .B(n313), .C(n308), .Z(n304) );
  GTECH_NOR2 U254 ( .A(b[5]), .B(a[5]), .Z(n308) );
  GTECH_NOR2 U255 ( .A(a[4]), .B(b[4]), .Z(n313) );
  GTECH_NAND2 U256 ( .A(b[5]), .B(a[5]), .Z(n306) );
  GTECH_AOI21 U257 ( .A(n361), .B(a[11]), .C(n385), .Z(n377) );
  GTECH_OA21 U258 ( .A(a[11]), .B(n361), .C(b[11]), .Z(n385) );
  GTECH_NAND2 U259 ( .A(n386), .B(n364), .Z(n361) );
  GTECH_NAND2 U260 ( .A(a[10]), .B(b[10]), .Z(n364) );
  GTECH_OAI21 U261 ( .A(a[10]), .B(b[10]), .C(n371), .Z(n386) );
  GTECH_OAI2N2 U262 ( .A(n287), .B(n284), .C(a[9]), .D(b[9]), .Z(n371) );
  GTECH_NOR2 U263 ( .A(b[8]), .B(a[8]), .Z(n284) );
  GTECH_NOR2 U264 ( .A(b[9]), .B(a[9]), .Z(n287) );
endmodule

