
module carry_select_adder8 ( a, b, cin, cout, sum );
  input [7:0] a;
  input [7:0] b;
  output [7:0] sum;
  input cin;
  output cout;
  wire   n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181;

  GTECH_MUX2 U64 ( .A(n133), .B(n134), .S(n135), .Z(sum[7]) );
  GTECH_ADD_AB U65 ( .A(n136), .B(n137), .S(n134) );
  GTECH_AOI21 U66 ( .A(n138), .B(n139), .C(n140), .Z(n136) );
  GTECH_XNOR2 U67 ( .A(n141), .B(n137), .Z(n133) );
  GTECH_XNOR2 U68 ( .A(b[7]), .B(a[7]), .Z(n137) );
  GTECH_MUX2 U69 ( .A(n142), .B(n143), .S(n135), .Z(sum[6]) );
  GTECH_XNOR2 U70 ( .A(n144), .B(n139), .Z(n143) );
  GTECH_OAI21 U71 ( .A(n145), .B(n146), .C(n147), .Z(n139) );
  GTECH_XNOR2 U72 ( .A(n144), .B(n148), .Z(n142) );
  GTECH_OR_NOT U73 ( .A(n140), .B(n138), .Z(n144) );
  GTECH_MUX2 U74 ( .A(n149), .B(n150), .S(n151), .Z(sum[5]) );
  GTECH_OA21 U75 ( .A(n152), .B(n135), .C(n146), .Z(n151) );
  GTECH_ADD_AB U76 ( .A(b[5]), .B(a[5]), .S(n150) );
  GTECH_OR_NOT U77 ( .A(n145), .B(n147), .Z(n149) );
  GTECH_OAI21 U78 ( .A(n153), .B(n135), .C(n154), .Z(sum[4]) );
  GTECH_MUX2 U79 ( .A(n155), .B(n156), .S(cin), .Z(sum[3]) );
  GTECH_ADD_AB U80 ( .A(n157), .B(n158), .S(n156) );
  GTECH_ADD_AB U81 ( .A(n159), .B(n158), .S(n155) );
  GTECH_ADD_AB U82 ( .A(b[3]), .B(a[3]), .S(n158) );
  GTECH_OA21 U83 ( .A(a[2]), .B(n160), .C(n161), .Z(n159) );
  GTECH_AO21 U84 ( .A(n160), .B(a[2]), .C(b[2]), .Z(n161) );
  GTECH_MUX2 U85 ( .A(n162), .B(n163), .S(cin), .Z(sum[2]) );
  GTECH_XNOR2 U86 ( .A(n164), .B(n165), .Z(n163) );
  GTECH_XNOR2 U87 ( .A(n160), .B(n165), .Z(n162) );
  GTECH_XNOR2 U88 ( .A(b[2]), .B(a[2]), .Z(n165) );
  GTECH_AO21 U89 ( .A(n166), .B(n167), .C(n168), .Z(n160) );
  GTECH_MUX2 U90 ( .A(n169), .B(n170), .S(n171), .Z(sum[1]) );
  GTECH_AND_NOT U91 ( .A(n166), .B(n168), .Z(n171) );
  GTECH_OAI21 U92 ( .A(cin), .B(n167), .C(n172), .Z(n170) );
  GTECH_AO21 U93 ( .A(n172), .B(cin), .C(n167), .Z(n169) );
  GTECH_AND2 U94 ( .A(b[0]), .B(a[0]), .Z(n167) );
  GTECH_ADD_AB U95 ( .A(cin), .B(n173), .S(sum[0]) );
  GTECH_OAI21 U96 ( .A(n174), .B(n135), .C(n154), .Z(cout) );
  GTECH_NAND2 U97 ( .A(n135), .B(n153), .Z(n154) );
  GTECH_AND_NOT U98 ( .A(n146), .B(n152), .Z(n153) );
  GTECH_NAND2 U99 ( .A(b[4]), .B(a[4]), .Z(n146) );
  GTECH_NOT U100 ( .A(n175), .Z(n135) );
  GTECH_MUX2 U101 ( .A(n173), .B(n176), .S(cin), .Z(n175) );
  GTECH_OA21 U102 ( .A(a[3]), .B(n157), .C(n177), .Z(n176) );
  GTECH_AO21 U103 ( .A(n157), .B(a[3]), .C(b[3]), .Z(n177) );
  GTECH_AO21 U104 ( .A(n164), .B(a[2]), .C(n178), .Z(n157) );
  GTECH_OA21 U105 ( .A(a[2]), .B(n164), .C(b[2]), .Z(n178) );
  GTECH_AO21 U106 ( .A(n166), .B(n172), .C(n168), .Z(n164) );
  GTECH_AND2 U107 ( .A(a[1]), .B(b[1]), .Z(n168) );
  GTECH_OR2 U108 ( .A(b[0]), .B(a[0]), .Z(n172) );
  GTECH_OR2 U109 ( .A(b[1]), .B(a[1]), .Z(n166) );
  GTECH_ADD_AB U110 ( .A(b[0]), .B(a[0]), .S(n173) );
  GTECH_AOI21 U111 ( .A(n141), .B(a[7]), .C(n179), .Z(n174) );
  GTECH_OA21 U112 ( .A(a[7]), .B(n141), .C(b[7]), .Z(n179) );
  GTECH_AO21 U113 ( .A(n138), .B(n148), .C(n140), .Z(n141) );
  GTECH_AND2 U114 ( .A(a[6]), .B(b[6]), .Z(n140) );
  GTECH_OAI21 U115 ( .A(n145), .B(n152), .C(n147), .Z(n148) );
  GTECH_NAND2 U116 ( .A(b[5]), .B(a[5]), .Z(n147) );
  GTECH_AND_NOT U117 ( .A(n180), .B(a[4]), .Z(n152) );
  GTECH_NOT U118 ( .A(b[4]), .Z(n180) );
  GTECH_AND_NOT U119 ( .A(n181), .B(a[5]), .Z(n145) );
  GTECH_NOT U120 ( .A(b[5]), .Z(n181) );
  GTECH_OR2 U121 ( .A(a[6]), .B(b[6]), .Z(n138) );
endmodule

