
module carry_ahead_adder16 ( a, b, cin, cout, sum, Gm, Pm );
  input [15:0] a;
  input [15:0] b;
  output [15:0] sum;
  input cin;
  output cout, Gm, Pm;
  wire   n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148;

  GTECH_ADD_AB U92 ( .A(n73), .B(n74), .S(sum[9]) );
  GTECH_ADD_AB U93 ( .A(n75), .B(n76), .S(sum[8]) );
  GTECH_ADD_AB U94 ( .A(n77), .B(n78), .S(sum[7]) );
  GTECH_OA21 U95 ( .A(n79), .B(n80), .C(n81), .Z(n78) );
  GTECH_ADD_AB U96 ( .A(n79), .B(n80), .S(sum[6]) );
  GTECH_OA21 U97 ( .A(n82), .B(n83), .C(n84), .Z(n79) );
  GTECH_ADD_AB U98 ( .A(n82), .B(n83), .S(sum[5]) );
  GTECH_OA21 U99 ( .A(n85), .B(n86), .C(n87), .Z(n82) );
  GTECH_ADD_AB U100 ( .A(n85), .B(n86), .S(sum[4]) );
  GTECH_XNOR2 U101 ( .A(n88), .B(n89), .Z(sum[3]) );
  GTECH_AOI21 U102 ( .A(n90), .B(n91), .C(n92), .Z(n88) );
  GTECH_ADD_AB U103 ( .A(n91), .B(n90), .S(sum[2]) );
  GTECH_AO21 U104 ( .A(n93), .B(n94), .C(n95), .Z(n90) );
  GTECH_ADD_AB U105 ( .A(n94), .B(n93), .S(sum[1]) );
  GTECH_AO21 U106 ( .A(n96), .B(cin), .C(n97), .Z(n93) );
  GTECH_ADD_AB U107 ( .A(n98), .B(n99), .S(sum[15]) );
  GTECH_AOI21 U108 ( .A(n100), .B(n101), .C(n102), .Z(n99) );
  GTECH_XNOR2 U109 ( .A(n100), .B(n103), .Z(sum[14]) );
  GTECH_OAI21 U110 ( .A(n104), .B(n105), .C(n106), .Z(n100) );
  GTECH_ADD_AB U111 ( .A(n104), .B(n105), .S(sum[13]) );
  GTECH_OA21 U112 ( .A(n107), .B(n108), .C(n109), .Z(n104) );
  GTECH_XNOR2 U113 ( .A(cout), .B(n108), .Z(sum[12]) );
  GTECH_ADD_AB U114 ( .A(n110), .B(n111), .S(sum[11]) );
  GTECH_AOI21 U115 ( .A(n112), .B(n113), .C(n114), .Z(n111) );
  GTECH_ADD_AB U116 ( .A(n113), .B(n112), .S(sum[10]) );
  GTECH_OAI21 U117 ( .A(n73), .B(n74), .C(n115), .Z(n112) );
  GTECH_OA21 U118 ( .A(n75), .B(n76), .C(n116), .Z(n73) );
  GTECH_ADD_AB U119 ( .A(cin), .B(n96), .S(sum[0]) );
  GTECH_NOT U120 ( .A(n107), .Z(cout) );
  GTECH_OA21 U121 ( .A(n75), .B(n117), .C(n118), .Z(n107) );
  GTECH_OA21 U122 ( .A(n85), .B(n119), .C(n120), .Z(n75) );
  GTECH_AND2 U123 ( .A(n121), .B(n122), .Z(n85) );
  GTECH_NAND4 U124 ( .A(n96), .B(n123), .C(cin), .D(n124), .Z(n121) );
  GTECH_AND3 U125 ( .A(n94), .B(n89), .C(n91), .Z(n124) );
  GTECH_AND4 U126 ( .A(n125), .B(n96), .C(n126), .D(n127), .Z(Pm) );
  GTECH_AND4 U127 ( .A(n123), .B(n91), .C(n94), .D(n89), .Z(n127) );
  GTECH_OA21 U128 ( .A(a[0]), .B(b[0]), .C(n128), .Z(n96) );
  GTECH_NOT U129 ( .A(n119), .Z(n125) );
  GTECH_OAI21 U130 ( .A(n129), .B(n117), .C(n118), .Z(Gm) );
  GTECH_OA21 U131 ( .A(n130), .B(n98), .C(n131), .Z(n118) );
  GTECH_AOI21 U132 ( .A(n132), .B(n101), .C(n102), .Z(n130) );
  GTECH_OAI21 U133 ( .A(n109), .B(n105), .C(n106), .Z(n132) );
  GTECH_NOT U134 ( .A(n126), .Z(n117) );
  GTECH_NOR4 U135 ( .A(n108), .B(n98), .C(n103), .D(n105), .Z(n126) );
  GTECH_OAI21 U136 ( .A(b[13]), .B(a[13]), .C(n106), .Z(n105) );
  GTECH_NAND2 U137 ( .A(b[13]), .B(a[13]), .Z(n106) );
  GTECH_NOT U138 ( .A(n101), .Z(n103) );
  GTECH_OA21 U139 ( .A(b[14]), .B(a[14]), .C(n133), .Z(n101) );
  GTECH_NOT U140 ( .A(n102), .Z(n133) );
  GTECH_AND2 U141 ( .A(b[14]), .B(a[14]), .Z(n102) );
  GTECH_OAI21 U142 ( .A(b[15]), .B(a[15]), .C(n131), .Z(n98) );
  GTECH_NAND2 U143 ( .A(a[15]), .B(b[15]), .Z(n131) );
  GTECH_OAI21 U144 ( .A(b[12]), .B(a[12]), .C(n109), .Z(n108) );
  GTECH_NAND2 U145 ( .A(a[12]), .B(b[12]), .Z(n109) );
  GTECH_OA21 U146 ( .A(n122), .B(n119), .C(n120), .Z(n129) );
  GTECH_OA21 U147 ( .A(n134), .B(n110), .C(n135), .Z(n120) );
  GTECH_AOI21 U148 ( .A(n136), .B(n113), .C(n114), .Z(n134) );
  GTECH_NOT U149 ( .A(n137), .Z(n113) );
  GTECH_OAI21 U150 ( .A(n116), .B(n74), .C(n115), .Z(n136) );
  GTECH_OR4 U151 ( .A(n76), .B(n110), .C(n137), .D(n74), .Z(n119) );
  GTECH_OAI21 U152 ( .A(b[9]), .B(a[9]), .C(n115), .Z(n74) );
  GTECH_NAND2 U153 ( .A(a[9]), .B(b[9]), .Z(n115) );
  GTECH_OAI21 U154 ( .A(b[10]), .B(a[10]), .C(n138), .Z(n137) );
  GTECH_NOT U155 ( .A(n114), .Z(n138) );
  GTECH_AND2 U156 ( .A(b[10]), .B(a[10]), .Z(n114) );
  GTECH_OAI21 U157 ( .A(b[11]), .B(a[11]), .C(n135), .Z(n110) );
  GTECH_NAND2 U158 ( .A(a[11]), .B(b[11]), .Z(n135) );
  GTECH_OAI21 U159 ( .A(b[8]), .B(a[8]), .C(n116), .Z(n76) );
  GTECH_NAND2 U160 ( .A(a[8]), .B(b[8]), .Z(n116) );
  GTECH_OA21 U161 ( .A(n139), .B(n140), .C(n141), .Z(n122) );
  GTECH_OA21 U162 ( .A(n142), .B(n77), .C(n143), .Z(n141) );
  GTECH_OA21 U163 ( .A(n144), .B(n80), .C(n81), .Z(n142) );
  GTECH_OA21 U164 ( .A(n83), .B(n87), .C(n84), .Z(n144) );
  GTECH_NOT U165 ( .A(n123), .Z(n140) );
  GTECH_NOR4 U166 ( .A(n86), .B(n77), .C(n80), .D(n83), .Z(n123) );
  GTECH_OAI21 U167 ( .A(b[5]), .B(a[5]), .C(n84), .Z(n83) );
  GTECH_NAND2 U168 ( .A(b[5]), .B(a[5]), .Z(n84) );
  GTECH_OAI21 U169 ( .A(b[6]), .B(a[6]), .C(n81), .Z(n80) );
  GTECH_NAND2 U170 ( .A(b[6]), .B(a[6]), .Z(n81) );
  GTECH_OAI21 U171 ( .A(b[7]), .B(a[7]), .C(n143), .Z(n77) );
  GTECH_NAND2 U172 ( .A(a[7]), .B(b[7]), .Z(n143) );
  GTECH_OAI21 U173 ( .A(b[4]), .B(a[4]), .C(n87), .Z(n86) );
  GTECH_NAND2 U174 ( .A(a[4]), .B(b[4]), .Z(n87) );
  GTECH_AOI22 U175 ( .A(b[3]), .B(a[3]), .C(n145), .D(n89), .Z(n139) );
  GTECH_ADD_AB U176 ( .A(b[3]), .B(a[3]), .S(n89) );
  GTECH_AO21 U177 ( .A(n146), .B(n91), .C(n92), .Z(n145) );
  GTECH_OA21 U178 ( .A(a[2]), .B(b[2]), .C(n147), .Z(n91) );
  GTECH_NOT U179 ( .A(n92), .Z(n147) );
  GTECH_AND2 U180 ( .A(b[2]), .B(a[2]), .Z(n92) );
  GTECH_AO21 U181 ( .A(n97), .B(n94), .C(n95), .Z(n146) );
  GTECH_NOT U182 ( .A(n148), .Z(n95) );
  GTECH_OA21 U183 ( .A(a[1]), .B(b[1]), .C(n148), .Z(n94) );
  GTECH_NAND2 U184 ( .A(a[1]), .B(b[1]), .Z(n148) );
  GTECH_NOT U185 ( .A(n128), .Z(n97) );
  GTECH_NAND2 U186 ( .A(a[0]), .B(b[0]), .Z(n128) );
endmodule

