
module booth_multiplier4 ( Rst, clk, Ld, M, R, Valid, P );
  input [15:0] M;
  input [15:0] R;
  output [31:0] P;
  input Rst, clk, Ld;
  output Valid;
  wire   N14, N15, N16, N17, N18, N19, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N41, N42, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N115, N116, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N155, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n127, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530;
  wire   [4:0] Cntr;
  wire   [16:0] A;
  wire   [33:0] Prod;

  GTECH_FJK1S Cntr_reg_0_ ( .J(n127), .K(n127), .TI(N14), .TE(N18), .CP(clk), 
        .Q(Cntr[0]), .QN(n264) );
  GTECH_FJK1S Cntr_reg_1_ ( .J(n127), .K(n127), .TI(N15), .TE(N18), .CP(clk), 
        .Q(Cntr[1]), .QN(n6) );
  GTECH_FJK1S Cntr_reg_2_ ( .J(n127), .K(n127), .TI(N16), .TE(N18), .CP(clk), 
        .Q(Cntr[2]), .QN(n7) );
  GTECH_FJK1S Cntr_reg_3_ ( .J(n127), .K(n127), .TI(N17), .TE(N18), .CP(clk), 
        .Q(Cntr[3]), .QN(n8) );
  GTECH_FJK1S Cntr_reg_4_ ( .J(n127), .K(n127), .TI(N19), .TE(N18), .CP(clk), 
        .Q(Cntr[4]), .QN(n9) );
  GTECH_FJK1S A_reg_16_ ( .J(n127), .K(n127), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[16]) );
  GTECH_FJK1S A_reg_15_ ( .J(n127), .K(n127), .TI(N42), .TE(N41), .CP(clk), 
        .Q(A[15]), .QN(n280) );
  GTECH_FJK1S A_reg_14_ ( .J(n127), .K(n127), .TI(N39), .TE(N41), .CP(clk), 
        .Q(A[14]), .QN(n279) );
  GTECH_FJK1S A_reg_13_ ( .J(n127), .K(n127), .TI(N38), .TE(N41), .CP(clk), 
        .Q(A[13]), .QN(n278) );
  GTECH_FJK1S A_reg_12_ ( .J(n127), .K(n127), .TI(N37), .TE(N41), .CP(clk), 
        .Q(A[12]), .QN(n277) );
  GTECH_FJK1S A_reg_11_ ( .J(n127), .K(n127), .TI(N36), .TE(N41), .CP(clk), 
        .Q(A[11]), .QN(n276) );
  GTECH_FJK1S A_reg_10_ ( .J(n127), .K(n127), .TI(N35), .TE(N41), .CP(clk), 
        .Q(A[10]), .QN(n275) );
  GTECH_FJK1S A_reg_9_ ( .J(n127), .K(n127), .TI(N34), .TE(N41), .CP(clk), .Q(
        A[9]), .QN(n274) );
  GTECH_FJK1S A_reg_8_ ( .J(n127), .K(n127), .TI(N33), .TE(N41), .CP(clk), .Q(
        A[8]), .QN(n273) );
  GTECH_FJK1S A_reg_7_ ( .J(n127), .K(n127), .TI(N32), .TE(N41), .CP(clk), .Q(
        A[7]), .QN(n272) );
  GTECH_FJK1S A_reg_6_ ( .J(n127), .K(n127), .TI(N31), .TE(N41), .CP(clk), .Q(
        A[6]), .QN(n271) );
  GTECH_FJK1S A_reg_5_ ( .J(n127), .K(n127), .TI(N30), .TE(N41), .CP(clk), .Q(
        A[5]), .QN(n270) );
  GTECH_FJK1S A_reg_4_ ( .J(n127), .K(n127), .TI(N29), .TE(N41), .CP(clk), .Q(
        A[4]), .QN(n269) );
  GTECH_FJK1S A_reg_3_ ( .J(n127), .K(n127), .TI(N28), .TE(N41), .CP(clk), .Q(
        A[3]), .QN(n268) );
  GTECH_FJK1S A_reg_2_ ( .J(n127), .K(n127), .TI(N27), .TE(N41), .CP(clk), .Q(
        A[2]), .QN(n267) );
  GTECH_FJK1S A_reg_1_ ( .J(n127), .K(n127), .TI(N26), .TE(N41), .CP(clk), .Q(
        A[1]), .QN(n266) );
  GTECH_FJK1S A_reg_0_ ( .J(n127), .K(n127), .TI(N25), .TE(N41), .CP(clk), .Q(
        A[0]), .QN(n265) );
  GTECH_FJK1S Prod_reg_0_ ( .J(n127), .K(n127), .TI(N82), .TE(N115), .CP(clk), 
        .Q(Prod[0]), .QN(n10) );
  GTECH_FJK1S Prod_reg_18_ ( .J(n127), .K(n127), .TI(N100), .TE(N115), .CP(clk), .Q(Prod[18]), .QN(n11) );
  GTECH_FJK1S Prod_reg_17_ ( .J(n127), .K(n127), .TI(N99), .TE(N115), .CP(clk), 
        .Q(Prod[17]), .QN(n12) );
  GTECH_FJK1S Prod_reg_16_ ( .J(n127), .K(n127), .TI(N98), .TE(N115), .CP(clk), 
        .Q(Prod[16]), .QN(n13) );
  GTECH_FJK1S Prod_reg_15_ ( .J(n127), .K(n127), .TI(N97), .TE(N115), .CP(clk), 
        .Q(Prod[15]), .QN(n14) );
  GTECH_FJK1S Prod_reg_14_ ( .J(n127), .K(n127), .TI(N96), .TE(N115), .CP(clk), 
        .Q(Prod[14]), .QN(n15) );
  GTECH_FJK1S Prod_reg_13_ ( .J(n127), .K(n127), .TI(N95), .TE(N115), .CP(clk), 
        .Q(Prod[13]), .QN(n16) );
  GTECH_FJK1S Prod_reg_12_ ( .J(n127), .K(n127), .TI(N94), .TE(N115), .CP(clk), 
        .Q(Prod[12]), .QN(n17) );
  GTECH_FJK1S Prod_reg_11_ ( .J(n127), .K(n127), .TI(N93), .TE(N115), .CP(clk), 
        .Q(Prod[11]), .QN(n18) );
  GTECH_FJK1S Prod_reg_10_ ( .J(n127), .K(n127), .TI(N92), .TE(N115), .CP(clk), 
        .Q(Prod[10]), .QN(n19) );
  GTECH_FJK1S Prod_reg_9_ ( .J(n127), .K(n127), .TI(N91), .TE(N115), .CP(clk), 
        .Q(Prod[9]), .QN(n20) );
  GTECH_FJK1S Prod_reg_8_ ( .J(n127), .K(n127), .TI(N90), .TE(N115), .CP(clk), 
        .Q(Prod[8]), .QN(n21) );
  GTECH_FJK1S Prod_reg_7_ ( .J(n127), .K(n127), .TI(N89), .TE(N115), .CP(clk), 
        .Q(Prod[7]), .QN(n22) );
  GTECH_FJK1S Prod_reg_6_ ( .J(n127), .K(n127), .TI(N88), .TE(N115), .CP(clk), 
        .Q(Prod[6]), .QN(n23) );
  GTECH_FJK1S Prod_reg_5_ ( .J(n127), .K(n127), .TI(N87), .TE(N115), .CP(clk), 
        .Q(Prod[5]), .QN(n24) );
  GTECH_FJK1S Prod_reg_4_ ( .J(n127), .K(n127), .TI(N86), .TE(N115), .CP(clk), 
        .Q(Prod[4]), .QN(n25) );
  GTECH_FJK1S Prod_reg_3_ ( .J(n127), .K(n127), .TI(N85), .TE(N115), .CP(clk), 
        .Q(Prod[3]), .QN(n26) );
  GTECH_FJK1S Prod_reg_2_ ( .J(n127), .K(n127), .TI(N84), .TE(N115), .CP(clk), 
        .Q(Prod[2]), .QN(n27) );
  GTECH_FJK1S Prod_reg_1_ ( .J(n127), .K(n127), .TI(N83), .TE(N115), .CP(clk), 
        .Q(Prod[1]), .QN(n28) );
  GTECH_FJK1S Prod_reg_19_ ( .J(n127), .K(n127), .TI(N101), .TE(N115), .CP(clk), .Q(Prod[19]), .QN(n29) );
  GTECH_FJK1S Prod_reg_33_ ( .J(n127), .K(n127), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[33]), .QN(n30) );
  GTECH_FJK1S Prod_reg_32_ ( .J(n127), .K(n127), .TI(N116), .TE(N115), .CP(clk), .Q(Prod[32]), .QN(n31) );
  GTECH_FJK1S Prod_reg_31_ ( .J(n127), .K(n127), .TI(N113), .TE(N115), .CP(clk), .Q(Prod[31]), .QN(n32) );
  GTECH_FJK1S Prod_reg_30_ ( .J(n127), .K(n127), .TI(N112), .TE(N115), .CP(clk), .Q(Prod[30]), .QN(n33) );
  GTECH_FJK1S Prod_reg_29_ ( .J(n127), .K(n127), .TI(N111), .TE(N115), .CP(clk), .Q(Prod[29]), .QN(n34) );
  GTECH_FJK1S Prod_reg_28_ ( .J(n127), .K(n127), .TI(N110), .TE(N115), .CP(clk), .Q(Prod[28]), .QN(n35) );
  GTECH_FJK1S Prod_reg_27_ ( .J(n127), .K(n127), .TI(N109), .TE(N115), .CP(clk), .Q(Prod[27]), .QN(n36) );
  GTECH_FJK1S Prod_reg_26_ ( .J(n127), .K(n127), .TI(N108), .TE(N115), .CP(clk), .Q(Prod[26]), .QN(n37) );
  GTECH_FJK1S Prod_reg_25_ ( .J(n127), .K(n127), .TI(N107), .TE(N115), .CP(clk), .Q(Prod[25]), .QN(n38) );
  GTECH_FJK1S Prod_reg_24_ ( .J(n127), .K(n127), .TI(N106), .TE(N115), .CP(clk), .Q(Prod[24]), .QN(n39) );
  GTECH_FJK1S Prod_reg_23_ ( .J(n127), .K(n127), .TI(N105), .TE(N115), .CP(clk), .Q(Prod[23]), .QN(n40) );
  GTECH_FJK1S Prod_reg_22_ ( .J(n127), .K(n127), .TI(N104), .TE(N115), .CP(clk), .Q(Prod[22]), .QN(n41) );
  GTECH_FJK1S Prod_reg_21_ ( .J(n127), .K(n127), .TI(N103), .TE(N115), .CP(clk), .Q(Prod[21]), .QN(n42) );
  GTECH_FJK1S Prod_reg_20_ ( .J(n127), .K(n127), .TI(N102), .TE(N115), .CP(clk), .Q(Prod[20]), .QN(n43) );
  GTECH_FJK1S P_reg_31_ ( .J(n127), .K(n127), .TI(N152), .TE(N151), .CP(clk), 
        .Q(P[31]) );
  GTECH_FJK1S P_reg_30_ ( .J(n127), .K(n127), .TI(N150), .TE(N151), .CP(clk), 
        .Q(P[30]) );
  GTECH_FJK1S P_reg_29_ ( .J(n127), .K(n127), .TI(N149), .TE(N151), .CP(clk), 
        .Q(P[29]) );
  GTECH_FJK1S P_reg_28_ ( .J(n127), .K(n127), .TI(N148), .TE(N151), .CP(clk), 
        .Q(P[28]) );
  GTECH_FJK1S P_reg_27_ ( .J(n127), .K(n127), .TI(N147), .TE(N151), .CP(clk), 
        .Q(P[27]) );
  GTECH_FJK1S P_reg_26_ ( .J(n127), .K(n127), .TI(N146), .TE(N151), .CP(clk), 
        .Q(P[26]) );
  GTECH_FJK1S P_reg_25_ ( .J(n127), .K(n127), .TI(N145), .TE(N151), .CP(clk), 
        .Q(P[25]) );
  GTECH_FJK1S P_reg_24_ ( .J(n127), .K(n127), .TI(N144), .TE(N151), .CP(clk), 
        .Q(P[24]) );
  GTECH_FJK1S P_reg_23_ ( .J(n127), .K(n127), .TI(N143), .TE(N151), .CP(clk), 
        .Q(P[23]) );
  GTECH_FJK1S P_reg_22_ ( .J(n127), .K(n127), .TI(N142), .TE(N151), .CP(clk), 
        .Q(P[22]) );
  GTECH_FJK1S P_reg_21_ ( .J(n127), .K(n127), .TI(N141), .TE(N151), .CP(clk), 
        .Q(P[21]) );
  GTECH_FJK1S P_reg_20_ ( .J(n127), .K(n127), .TI(N140), .TE(N151), .CP(clk), 
        .Q(P[20]) );
  GTECH_FJK1S P_reg_19_ ( .J(n127), .K(n127), .TI(N139), .TE(N151), .CP(clk), 
        .Q(P[19]) );
  GTECH_FJK1S P_reg_18_ ( .J(n127), .K(n127), .TI(N138), .TE(N151), .CP(clk), 
        .Q(P[18]) );
  GTECH_FJK1S P_reg_17_ ( .J(n127), .K(n127), .TI(N137), .TE(N151), .CP(clk), 
        .Q(P[17]) );
  GTECH_FJK1S P_reg_16_ ( .J(n127), .K(n127), .TI(N136), .TE(N151), .CP(clk), 
        .Q(P[16]) );
  GTECH_FJK1S P_reg_15_ ( .J(n127), .K(n127), .TI(N135), .TE(N151), .CP(clk), 
        .Q(P[15]) );
  GTECH_FJK1S P_reg_14_ ( .J(n127), .K(n127), .TI(N134), .TE(N151), .CP(clk), 
        .Q(P[14]) );
  GTECH_FJK1S P_reg_13_ ( .J(n127), .K(n127), .TI(N133), .TE(N151), .CP(clk), 
        .Q(P[13]) );
  GTECH_FJK1S P_reg_12_ ( .J(n127), .K(n127), .TI(N132), .TE(N151), .CP(clk), 
        .Q(P[12]) );
  GTECH_FJK1S P_reg_11_ ( .J(n127), .K(n127), .TI(N131), .TE(N151), .CP(clk), 
        .Q(P[11]) );
  GTECH_FJK1S P_reg_10_ ( .J(n127), .K(n127), .TI(N130), .TE(N151), .CP(clk), 
        .Q(P[10]) );
  GTECH_FJK1S P_reg_9_ ( .J(n127), .K(n127), .TI(N129), .TE(N151), .CP(clk), 
        .Q(P[9]) );
  GTECH_FJK1S P_reg_8_ ( .J(n127), .K(n127), .TI(N128), .TE(N151), .CP(clk), 
        .Q(P[8]) );
  GTECH_FJK1S P_reg_7_ ( .J(n127), .K(n127), .TI(N127), .TE(N151), .CP(clk), 
        .Q(P[7]) );
  GTECH_FJK1S P_reg_6_ ( .J(n127), .K(n127), .TI(N126), .TE(N151), .CP(clk), 
        .Q(P[6]) );
  GTECH_FJK1S P_reg_5_ ( .J(n127), .K(n127), .TI(N125), .TE(N151), .CP(clk), 
        .Q(P[5]) );
  GTECH_FJK1S P_reg_4_ ( .J(n127), .K(n127), .TI(N124), .TE(N151), .CP(clk), 
        .Q(P[4]) );
  GTECH_FJK1S P_reg_3_ ( .J(n127), .K(n127), .TI(N123), .TE(N151), .CP(clk), 
        .Q(P[3]) );
  GTECH_FJK1S P_reg_2_ ( .J(n127), .K(n127), .TI(N122), .TE(N151), .CP(clk), 
        .Q(P[2]) );
  GTECH_FJK1S P_reg_1_ ( .J(n127), .K(n127), .TI(N121), .TE(N151), .CP(clk), 
        .Q(P[1]) );
  GTECH_FJK1S P_reg_0_ ( .J(n127), .K(n127), .TI(N120), .TE(N151), .CP(clk), 
        .Q(P[0]) );
  GTECH_FD1 Valid_reg ( .D(N155), .CP(clk), .Q(Valid) );
  GTECH_ZERO U266 ( .Z(n127) );
  GTECH_NOT U267 ( .A(n282), .Z(N99) );
  GTECH_AOI222 U268 ( .A(n283), .B(n284), .C(n285), .D(n286), .E(n287), .F(
        n288), .Z(n282) );
  GTECH_NOT U269 ( .A(n289), .Z(N98) );
  GTECH_AOI222 U270 ( .A(n285), .B(n290), .C(n291), .D(n292), .E(R[15]), .F(
        n293), .Z(n289) );
  GTECH_NAND2 U271 ( .A(n294), .B(n295), .Z(n291) );
  GTECH_AO22 U272 ( .A(n296), .B(n297), .C(R[14]), .D(n293), .Z(N97) );
  GTECH_AO22 U273 ( .A(n296), .B(n298), .C(R[13]), .D(n293), .Z(N96) );
  GTECH_AO22 U274 ( .A(n296), .B(n299), .C(R[12]), .D(n293), .Z(N95) );
  GTECH_AO22 U275 ( .A(n296), .B(n300), .C(R[11]), .D(n293), .Z(N94) );
  GTECH_AO22 U276 ( .A(n296), .B(n301), .C(R[10]), .D(n293), .Z(N93) );
  GTECH_AO22 U277 ( .A(n296), .B(n302), .C(R[9]), .D(n293), .Z(N92) );
  GTECH_AO22 U278 ( .A(n296), .B(n303), .C(R[8]), .D(n293), .Z(N91) );
  GTECH_AO22 U279 ( .A(n296), .B(n304), .C(R[7]), .D(n293), .Z(N90) );
  GTECH_AO22 U280 ( .A(n296), .B(n305), .C(R[6]), .D(n293), .Z(N89) );
  GTECH_AO22 U281 ( .A(n296), .B(n306), .C(R[5]), .D(n293), .Z(N88) );
  GTECH_AO22 U282 ( .A(n296), .B(n307), .C(R[4]), .D(n293), .Z(N87) );
  GTECH_AO22 U283 ( .A(n296), .B(n308), .C(R[3]), .D(n293), .Z(N86) );
  GTECH_AO22 U284 ( .A(n296), .B(n309), .C(R[2]), .D(n293), .Z(N85) );
  GTECH_AO22 U285 ( .A(n296), .B(n310), .C(R[1]), .D(n293), .Z(N84) );
  GTECH_AO22 U286 ( .A(n296), .B(n311), .C(R[0]), .D(n293), .Z(N83) );
  GTECH_AND2 U287 ( .A(M[15]), .B(n293), .Z(N42) );
  GTECH_AND2 U288 ( .A(M[14]), .B(n293), .Z(N39) );
  GTECH_AND2 U289 ( .A(M[13]), .B(n293), .Z(N38) );
  GTECH_AND2 U290 ( .A(M[12]), .B(n293), .Z(N37) );
  GTECH_AND2 U291 ( .A(M[11]), .B(n293), .Z(N36) );
  GTECH_AND2 U292 ( .A(M[10]), .B(n293), .Z(N35) );
  GTECH_AND2 U293 ( .A(M[9]), .B(n293), .Z(N34) );
  GTECH_AND2 U294 ( .A(M[8]), .B(n293), .Z(N33) );
  GTECH_AND2 U295 ( .A(M[7]), .B(n293), .Z(N32) );
  GTECH_AND2 U296 ( .A(M[6]), .B(n293), .Z(N31) );
  GTECH_AND2 U297 ( .A(M[5]), .B(n293), .Z(N30) );
  GTECH_AND2 U298 ( .A(M[4]), .B(n293), .Z(N29) );
  GTECH_AND2 U299 ( .A(M[3]), .B(n293), .Z(N28) );
  GTECH_AND2 U300 ( .A(M[2]), .B(n293), .Z(N27) );
  GTECH_AND2 U301 ( .A(M[1]), .B(n293), .Z(N26) );
  GTECH_AND2 U302 ( .A(M[0]), .B(n293), .Z(N25) );
  GTECH_NOT U303 ( .A(n312), .Z(n293) );
  GTECH_NAND2 U304 ( .A(n312), .B(n313), .Z(N19) );
  GTECH_NAND3 U305 ( .A(n314), .B(n315), .C(n296), .Z(n313) );
  GTECH_NAND3 U306 ( .A(n316), .B(n317), .C(n318), .Z(N18) );
  GTECH_AND2 U307 ( .A(n296), .B(n319), .Z(N17) );
  GTECH_OAI21 U308 ( .A(n8), .B(n320), .C(n314), .Z(n319) );
  GTECH_AND2 U309 ( .A(n296), .B(n321), .Z(N16) );
  GTECH_OAI21 U310 ( .A(n7), .B(n322), .C(n323), .Z(n321) );
  GTECH_NOT U311 ( .A(n324), .Z(N152) );
  GTECH_AOI222 U312 ( .A(n325), .B(n326), .C(n327), .D(n328), .E(n329), .F(
        n330), .Z(n324) );
  GTECH_NAND2 U313 ( .A(n317), .B(n331), .Z(N151) );
  GTECH_NOT U314 ( .A(n332), .Z(N150) );
  GTECH_AOI222 U315 ( .A(n333), .B(n325), .C(n327), .D(n334), .E(n329), .F(
        n335), .Z(n332) );
  GTECH_MUX2 U316 ( .A(n336), .B(N14), .S(n6), .Z(N15) );
  GTECH_AND_NOT U317 ( .A(n296), .B(n264), .Z(n336) );
  GTECH_NOT U318 ( .A(n337), .Z(N149) );
  GTECH_AOI222 U319 ( .A(n338), .B(n325), .C(n327), .D(n339), .E(n329), .F(
        n340), .Z(n337) );
  GTECH_NOT U320 ( .A(n341), .Z(N148) );
  GTECH_AOI222 U321 ( .A(n342), .B(n325), .C(n327), .D(n343), .E(n329), .F(
        n344), .Z(n341) );
  GTECH_NOT U322 ( .A(n345), .Z(N147) );
  GTECH_AOI222 U323 ( .A(n346), .B(n325), .C(n327), .D(n347), .E(n329), .F(
        n348), .Z(n345) );
  GTECH_NOT U324 ( .A(n349), .Z(N146) );
  GTECH_AOI222 U325 ( .A(n350), .B(n325), .C(n327), .D(n351), .E(n329), .F(
        n352), .Z(n349) );
  GTECH_NOT U326 ( .A(n353), .Z(N145) );
  GTECH_AOI222 U327 ( .A(n354), .B(n325), .C(n327), .D(n355), .E(n329), .F(
        n356), .Z(n353) );
  GTECH_NOT U328 ( .A(n357), .Z(N144) );
  GTECH_AOI222 U329 ( .A(n358), .B(n325), .C(n327), .D(n359), .E(n329), .F(
        n360), .Z(n357) );
  GTECH_NOT U330 ( .A(n361), .Z(N143) );
  GTECH_AOI222 U331 ( .A(n362), .B(n325), .C(n327), .D(n363), .E(n329), .F(
        n364), .Z(n361) );
  GTECH_NOT U332 ( .A(n365), .Z(N142) );
  GTECH_AOI222 U333 ( .A(n366), .B(n325), .C(n327), .D(n367), .E(n329), .F(
        n368), .Z(n365) );
  GTECH_NOT U334 ( .A(n369), .Z(N141) );
  GTECH_AOI222 U335 ( .A(n370), .B(n325), .C(n327), .D(n371), .E(n329), .F(
        n372), .Z(n369) );
  GTECH_NOT U336 ( .A(n373), .Z(N140) );
  GTECH_AOI222 U337 ( .A(n374), .B(n325), .C(n327), .D(n375), .E(n329), .F(
        n376), .Z(n373) );
  GTECH_NOT U338 ( .A(n377), .Z(N14) );
  GTECH_NAND2 U339 ( .A(n296), .B(n264), .Z(n377) );
  GTECH_NOT U340 ( .A(n378), .Z(N139) );
  GTECH_AOI222 U341 ( .A(n379), .B(n325), .C(n327), .D(n380), .E(n329), .F(
        n381), .Z(n378) );
  GTECH_NOT U342 ( .A(n382), .Z(N138) );
  GTECH_AOI222 U343 ( .A(n383), .B(n325), .C(n327), .D(n384), .E(n329), .F(
        n385), .Z(n382) );
  GTECH_NOT U344 ( .A(n386), .Z(N137) );
  GTECH_AOI222 U345 ( .A(n387), .B(n325), .C(n327), .D(n388), .E(n329), .F(
        n389), .Z(n386) );
  GTECH_NOT U346 ( .A(n390), .Z(N136) );
  GTECH_AOI222 U347 ( .A(n325), .B(n284), .C(n327), .D(n286), .E(n329), .F(
        n288), .Z(n390) );
  GTECH_NOT U348 ( .A(n391), .Z(n288) );
  GTECH_XOR2 U349 ( .A(n392), .B(n393), .Z(n391) );
  GTECH_NOT U350 ( .A(n394), .Z(n393) );
  GTECH_NOT U351 ( .A(n395), .Z(n327) );
  GTECH_NOT U352 ( .A(n396), .Z(n284) );
  GTECH_XOR2 U353 ( .A(n392), .B(n397), .Z(n396) );
  GTECH_NOT U354 ( .A(n398), .Z(n397) );
  GTECH_XOR2 U355 ( .A(n286), .B(n266), .Z(n392) );
  GTECH_OAI21 U356 ( .A(n12), .B(n395), .C(n399), .Z(N135) );
  GTECH_OAI21 U357 ( .A(n329), .B(n325), .C(n292), .Z(n399) );
  GTECH_OAI21 U358 ( .A(n12), .B(n400), .C(n394), .Z(n292) );
  GTECH_NOT U359 ( .A(n401), .Z(n325) );
  GTECH_NAND3 U360 ( .A(n28), .B(n402), .C(N155), .Z(n401) );
  GTECH_NOT U361 ( .A(n403), .Z(n329) );
  GTECH_NAND3 U362 ( .A(n10), .B(n404), .C(N155), .Z(n403) );
  GTECH_NAND2 U363 ( .A(n405), .B(N155), .Z(n395) );
  GTECH_XOR2 U364 ( .A(n402), .B(n28), .Z(n405) );
  GTECH_AND2 U365 ( .A(N155), .B(n297), .Z(N134) );
  GTECH_NOT U366 ( .A(n13), .Z(n297) );
  GTECH_AND2 U367 ( .A(N155), .B(n298), .Z(N133) );
  GTECH_NOT U368 ( .A(n14), .Z(n298) );
  GTECH_AND2 U369 ( .A(N155), .B(n299), .Z(N132) );
  GTECH_NOT U370 ( .A(n15), .Z(n299) );
  GTECH_AND2 U371 ( .A(N155), .B(n300), .Z(N131) );
  GTECH_NOT U372 ( .A(n16), .Z(n300) );
  GTECH_AND2 U373 ( .A(N155), .B(n301), .Z(N130) );
  GTECH_NOT U374 ( .A(n17), .Z(n301) );
  GTECH_AND2 U375 ( .A(N155), .B(n302), .Z(N129) );
  GTECH_NOT U376 ( .A(n18), .Z(n302) );
  GTECH_AND2 U377 ( .A(N155), .B(n303), .Z(N128) );
  GTECH_NOT U378 ( .A(n19), .Z(n303) );
  GTECH_AND2 U379 ( .A(N155), .B(n304), .Z(N127) );
  GTECH_NOT U380 ( .A(n20), .Z(n304) );
  GTECH_AND2 U381 ( .A(N155), .B(n305), .Z(N126) );
  GTECH_NOT U382 ( .A(n21), .Z(n305) );
  GTECH_AND2 U383 ( .A(N155), .B(n306), .Z(N125) );
  GTECH_NOT U384 ( .A(n22), .Z(n306) );
  GTECH_AND2 U385 ( .A(N155), .B(n307), .Z(N124) );
  GTECH_NOT U386 ( .A(n23), .Z(n307) );
  GTECH_AND2 U387 ( .A(N155), .B(n308), .Z(N123) );
  GTECH_NOT U388 ( .A(n24), .Z(n308) );
  GTECH_AND2 U389 ( .A(N155), .B(n309), .Z(N122) );
  GTECH_NOT U390 ( .A(n25), .Z(n309) );
  GTECH_AND2 U391 ( .A(N155), .B(n310), .Z(N121) );
  GTECH_NOT U392 ( .A(n26), .Z(n310) );
  GTECH_AND2 U393 ( .A(N155), .B(n311), .Z(N120) );
  GTECH_NOT U394 ( .A(n27), .Z(n311) );
  GTECH_NOT U395 ( .A(n331), .Z(N155) );
  GTECH_NAND5 U396 ( .A(n406), .B(n6), .C(n9), .D(n8), .E(n7), .Z(n331) );
  GTECH_NOR2 U397 ( .A(n264), .B(Rst), .Z(n406) );
  GTECH_NOT U398 ( .A(n407), .Z(N116) );
  GTECH_AOI222 U399 ( .A(n285), .B(n328), .C(n287), .D(n330), .E(n326), .F(
        n283), .Z(n407) );
  GTECH_XOR2 U400 ( .A(n408), .B(n409), .Z(n326) );
  GTECH_ADD_ABC U401 ( .A(n31), .B(n280), .C(n410), .COUT(n409) );
  GTECH_XOR2 U402 ( .A(n411), .B(n408), .Z(n330) );
  GTECH_XOR2 U403 ( .A(A[16]), .B(n30), .Z(n408) );
  GTECH_OAI21 U404 ( .A(n412), .B(n31), .C(n413), .Z(n411) );
  GTECH_OAI21 U405 ( .A(n280), .B(n334), .C(n414), .Z(n413) );
  GTECH_NOT U406 ( .A(n30), .Z(n328) );
  GTECH_NAND2 U407 ( .A(n318), .B(n415), .Z(N115) );
  GTECH_NOT U408 ( .A(N41), .Z(n415) );
  GTECH_NAND2 U409 ( .A(n317), .B(n312), .Z(N41) );
  GTECH_NAND2 U410 ( .A(Ld), .B(n317), .Z(n312) );
  GTECH_NOT U411 ( .A(n416), .Z(N113) );
  GTECH_AOI222 U412 ( .A(n285), .B(n334), .C(n287), .D(n335), .E(n333), .F(
        n283), .Z(n416) );
  GTECH_XOR2 U413 ( .A(n417), .B(n410), .Z(n333) );
  GTECH_ADD_ABC U414 ( .A(n32), .B(n279), .C(n418), .COUT(n410) );
  GTECH_NOT U415 ( .A(n419), .Z(n335) );
  GTECH_XOR2 U416 ( .A(n417), .B(n420), .Z(n419) );
  GTECH_NOT U417 ( .A(n414), .Z(n420) );
  GTECH_OAI21 U418 ( .A(n32), .B(n421), .C(n422), .Z(n414) );
  GTECH_OAI21 U419 ( .A(n279), .B(n339), .C(n423), .Z(n422) );
  GTECH_XOR2 U420 ( .A(n412), .B(n31), .Z(n417) );
  GTECH_NOT U421 ( .A(n280), .Z(n412) );
  GTECH_NOT U422 ( .A(n31), .Z(n334) );
  GTECH_NOT U423 ( .A(n424), .Z(N112) );
  GTECH_AOI222 U424 ( .A(n285), .B(n339), .C(n287), .D(n340), .E(n338), .F(
        n283), .Z(n424) );
  GTECH_XOR2 U425 ( .A(n425), .B(n418), .Z(n338) );
  GTECH_ADD_ABC U426 ( .A(n33), .B(n278), .C(n426), .COUT(n418) );
  GTECH_NOT U427 ( .A(n427), .Z(n340) );
  GTECH_XOR2 U428 ( .A(n425), .B(n428), .Z(n427) );
  GTECH_NOT U429 ( .A(n423), .Z(n428) );
  GTECH_OAI21 U430 ( .A(n33), .B(n429), .C(n430), .Z(n423) );
  GTECH_OAI21 U431 ( .A(n278), .B(n343), .C(n431), .Z(n430) );
  GTECH_XOR2 U432 ( .A(n421), .B(n32), .Z(n425) );
  GTECH_NOT U433 ( .A(n279), .Z(n421) );
  GTECH_NOT U434 ( .A(n32), .Z(n339) );
  GTECH_NOT U435 ( .A(n432), .Z(N111) );
  GTECH_AOI222 U436 ( .A(n285), .B(n343), .C(n287), .D(n344), .E(n342), .F(
        n283), .Z(n432) );
  GTECH_XOR2 U437 ( .A(n433), .B(n426), .Z(n342) );
  GTECH_ADD_ABC U438 ( .A(n34), .B(n277), .C(n434), .COUT(n426) );
  GTECH_NOT U439 ( .A(n435), .Z(n344) );
  GTECH_XOR2 U440 ( .A(n433), .B(n436), .Z(n435) );
  GTECH_NOT U441 ( .A(n431), .Z(n436) );
  GTECH_OAI21 U442 ( .A(n34), .B(n437), .C(n438), .Z(n431) );
  GTECH_OAI21 U443 ( .A(n277), .B(n347), .C(n439), .Z(n438) );
  GTECH_XOR2 U444 ( .A(n429), .B(n33), .Z(n433) );
  GTECH_NOT U445 ( .A(n278), .Z(n429) );
  GTECH_NOT U446 ( .A(n33), .Z(n343) );
  GTECH_NOT U447 ( .A(n440), .Z(N110) );
  GTECH_AOI222 U448 ( .A(n285), .B(n347), .C(n287), .D(n348), .E(n346), .F(
        n283), .Z(n440) );
  GTECH_XOR2 U449 ( .A(n441), .B(n434), .Z(n346) );
  GTECH_ADD_ABC U450 ( .A(n35), .B(n276), .C(n442), .COUT(n434) );
  GTECH_NOT U451 ( .A(n443), .Z(n348) );
  GTECH_XOR2 U452 ( .A(n441), .B(n444), .Z(n443) );
  GTECH_NOT U453 ( .A(n439), .Z(n444) );
  GTECH_OAI21 U454 ( .A(n35), .B(n445), .C(n446), .Z(n439) );
  GTECH_OAI21 U455 ( .A(n276), .B(n351), .C(n447), .Z(n446) );
  GTECH_XOR2 U456 ( .A(n437), .B(n34), .Z(n441) );
  GTECH_NOT U457 ( .A(n277), .Z(n437) );
  GTECH_NOT U458 ( .A(n34), .Z(n347) );
  GTECH_NOT U459 ( .A(n448), .Z(N109) );
  GTECH_AOI222 U460 ( .A(n285), .B(n351), .C(n287), .D(n352), .E(n350), .F(
        n283), .Z(n448) );
  GTECH_XOR2 U461 ( .A(n449), .B(n442), .Z(n350) );
  GTECH_ADD_ABC U462 ( .A(n36), .B(n275), .C(n450), .COUT(n442) );
  GTECH_NOT U463 ( .A(n451), .Z(n352) );
  GTECH_XOR2 U464 ( .A(n449), .B(n452), .Z(n451) );
  GTECH_NOT U465 ( .A(n447), .Z(n452) );
  GTECH_OAI21 U466 ( .A(n36), .B(n453), .C(n454), .Z(n447) );
  GTECH_OAI21 U467 ( .A(n275), .B(n355), .C(n455), .Z(n454) );
  GTECH_XOR2 U468 ( .A(n445), .B(n35), .Z(n449) );
  GTECH_NOT U469 ( .A(n276), .Z(n445) );
  GTECH_NOT U470 ( .A(n35), .Z(n351) );
  GTECH_NOT U471 ( .A(n456), .Z(N108) );
  GTECH_AOI222 U472 ( .A(n285), .B(n355), .C(n287), .D(n356), .E(n354), .F(
        n283), .Z(n456) );
  GTECH_XOR2 U473 ( .A(n457), .B(n450), .Z(n354) );
  GTECH_ADD_ABC U474 ( .A(n37), .B(n274), .C(n458), .COUT(n450) );
  GTECH_NOT U475 ( .A(n459), .Z(n356) );
  GTECH_XOR2 U476 ( .A(n457), .B(n460), .Z(n459) );
  GTECH_NOT U477 ( .A(n455), .Z(n460) );
  GTECH_OAI21 U478 ( .A(n37), .B(n461), .C(n462), .Z(n455) );
  GTECH_OAI21 U479 ( .A(n274), .B(n359), .C(n463), .Z(n462) );
  GTECH_XOR2 U480 ( .A(n453), .B(n36), .Z(n457) );
  GTECH_NOT U481 ( .A(n275), .Z(n453) );
  GTECH_NOT U482 ( .A(n36), .Z(n355) );
  GTECH_NOT U483 ( .A(n464), .Z(N107) );
  GTECH_AOI222 U484 ( .A(n285), .B(n359), .C(n287), .D(n360), .E(n358), .F(
        n283), .Z(n464) );
  GTECH_XOR2 U485 ( .A(n465), .B(n458), .Z(n358) );
  GTECH_ADD_ABC U486 ( .A(n38), .B(n273), .C(n466), .COUT(n458) );
  GTECH_NOT U487 ( .A(n467), .Z(n360) );
  GTECH_XOR2 U488 ( .A(n465), .B(n468), .Z(n467) );
  GTECH_NOT U489 ( .A(n463), .Z(n468) );
  GTECH_OAI21 U490 ( .A(n38), .B(n469), .C(n470), .Z(n463) );
  GTECH_OAI21 U491 ( .A(n273), .B(n363), .C(n471), .Z(n470) );
  GTECH_XOR2 U492 ( .A(n461), .B(n37), .Z(n465) );
  GTECH_NOT U493 ( .A(n274), .Z(n461) );
  GTECH_NOT U494 ( .A(n37), .Z(n359) );
  GTECH_NOT U495 ( .A(n472), .Z(N106) );
  GTECH_AOI222 U496 ( .A(n285), .B(n363), .C(n287), .D(n364), .E(n362), .F(
        n283), .Z(n472) );
  GTECH_XOR2 U497 ( .A(n473), .B(n466), .Z(n362) );
  GTECH_ADD_ABC U498 ( .A(n39), .B(n272), .C(n474), .COUT(n466) );
  GTECH_NOT U499 ( .A(n475), .Z(n364) );
  GTECH_XOR2 U500 ( .A(n473), .B(n476), .Z(n475) );
  GTECH_NOT U501 ( .A(n471), .Z(n476) );
  GTECH_OAI21 U502 ( .A(n39), .B(n477), .C(n478), .Z(n471) );
  GTECH_OAI21 U503 ( .A(n272), .B(n367), .C(n479), .Z(n478) );
  GTECH_XOR2 U504 ( .A(n469), .B(n38), .Z(n473) );
  GTECH_NOT U505 ( .A(n273), .Z(n469) );
  GTECH_NOT U506 ( .A(n38), .Z(n363) );
  GTECH_NOT U507 ( .A(n480), .Z(N105) );
  GTECH_AOI222 U508 ( .A(n285), .B(n367), .C(n287), .D(n368), .E(n366), .F(
        n283), .Z(n480) );
  GTECH_XOR2 U509 ( .A(n481), .B(n474), .Z(n366) );
  GTECH_ADD_ABC U510 ( .A(n40), .B(n271), .C(n482), .COUT(n474) );
  GTECH_NOT U511 ( .A(n483), .Z(n368) );
  GTECH_XOR2 U512 ( .A(n481), .B(n484), .Z(n483) );
  GTECH_NOT U513 ( .A(n479), .Z(n484) );
  GTECH_OAI21 U514 ( .A(n40), .B(n485), .C(n486), .Z(n479) );
  GTECH_OAI21 U515 ( .A(n271), .B(n371), .C(n487), .Z(n486) );
  GTECH_XOR2 U516 ( .A(n477), .B(n39), .Z(n481) );
  GTECH_NOT U517 ( .A(n272), .Z(n477) );
  GTECH_NOT U518 ( .A(n39), .Z(n367) );
  GTECH_NOT U519 ( .A(n488), .Z(N104) );
  GTECH_AOI222 U520 ( .A(n285), .B(n371), .C(n287), .D(n372), .E(n370), .F(
        n283), .Z(n488) );
  GTECH_XOR2 U521 ( .A(n489), .B(n482), .Z(n370) );
  GTECH_ADD_ABC U522 ( .A(n41), .B(n270), .C(n490), .COUT(n482) );
  GTECH_NOT U523 ( .A(n491), .Z(n372) );
  GTECH_XOR2 U524 ( .A(n489), .B(n492), .Z(n491) );
  GTECH_NOT U525 ( .A(n487), .Z(n492) );
  GTECH_OAI21 U526 ( .A(n41), .B(n493), .C(n494), .Z(n487) );
  GTECH_OAI21 U527 ( .A(n270), .B(n375), .C(n495), .Z(n494) );
  GTECH_XOR2 U528 ( .A(n485), .B(n40), .Z(n489) );
  GTECH_NOT U529 ( .A(n271), .Z(n485) );
  GTECH_NOT U530 ( .A(n40), .Z(n371) );
  GTECH_NOT U531 ( .A(n496), .Z(N103) );
  GTECH_AOI222 U532 ( .A(n285), .B(n375), .C(n287), .D(n376), .E(n374), .F(
        n283), .Z(n496) );
  GTECH_XOR2 U533 ( .A(n497), .B(n490), .Z(n374) );
  GTECH_ADD_ABC U534 ( .A(n42), .B(n269), .C(n498), .COUT(n490) );
  GTECH_NOT U535 ( .A(n499), .Z(n376) );
  GTECH_XOR2 U536 ( .A(n497), .B(n500), .Z(n499) );
  GTECH_NOT U537 ( .A(n495), .Z(n500) );
  GTECH_OAI21 U538 ( .A(n42), .B(n501), .C(n502), .Z(n495) );
  GTECH_OAI21 U539 ( .A(n269), .B(n380), .C(n503), .Z(n502) );
  GTECH_XOR2 U540 ( .A(n493), .B(n41), .Z(n497) );
  GTECH_NOT U541 ( .A(n270), .Z(n493) );
  GTECH_NOT U542 ( .A(n41), .Z(n375) );
  GTECH_NOT U543 ( .A(n504), .Z(N102) );
  GTECH_AOI222 U544 ( .A(n285), .B(n380), .C(n287), .D(n381), .E(n379), .F(
        n283), .Z(n504) );
  GTECH_XOR2 U545 ( .A(n505), .B(n498), .Z(n379) );
  GTECH_ADD_ABC U546 ( .A(n43), .B(n268), .C(n506), .COUT(n498) );
  GTECH_NOT U547 ( .A(n507), .Z(n381) );
  GTECH_XOR2 U548 ( .A(n505), .B(n508), .Z(n507) );
  GTECH_NOT U549 ( .A(n503), .Z(n508) );
  GTECH_OAI21 U550 ( .A(n43), .B(n509), .C(n510), .Z(n503) );
  GTECH_OAI21 U551 ( .A(n268), .B(n384), .C(n511), .Z(n510) );
  GTECH_XOR2 U552 ( .A(n501), .B(n42), .Z(n505) );
  GTECH_NOT U553 ( .A(n269), .Z(n501) );
  GTECH_NOT U554 ( .A(n42), .Z(n380) );
  GTECH_NOT U555 ( .A(n512), .Z(N101) );
  GTECH_AOI222 U556 ( .A(n285), .B(n384), .C(n287), .D(n385), .E(n383), .F(
        n283), .Z(n512) );
  GTECH_XOR2 U557 ( .A(n513), .B(n506), .Z(n383) );
  GTECH_ADD_ABC U558 ( .A(n29), .B(n267), .C(n514), .COUT(n506) );
  GTECH_NOT U559 ( .A(n515), .Z(n385) );
  GTECH_XOR2 U560 ( .A(n513), .B(n516), .Z(n515) );
  GTECH_NOT U561 ( .A(n511), .Z(n516) );
  GTECH_OAI21 U562 ( .A(n29), .B(n517), .C(n518), .Z(n511) );
  GTECH_OAI21 U563 ( .A(n267), .B(n388), .C(n519), .Z(n518) );
  GTECH_XOR2 U564 ( .A(n509), .B(n43), .Z(n513) );
  GTECH_NOT U565 ( .A(n268), .Z(n509) );
  GTECH_NOT U566 ( .A(n43), .Z(n384) );
  GTECH_NOT U567 ( .A(n520), .Z(N100) );
  GTECH_AOI222 U568 ( .A(n387), .B(n283), .C(n285), .D(n388), .E(n287), .F(
        n389), .Z(n520) );
  GTECH_NOT U569 ( .A(n521), .Z(n389) );
  GTECH_XOR2 U570 ( .A(n522), .B(n523), .Z(n521) );
  GTECH_NOT U571 ( .A(n519), .Z(n523) );
  GTECH_OAI21 U572 ( .A(n11), .B(n524), .C(n525), .Z(n519) );
  GTECH_OAI21 U573 ( .A(n266), .B(n286), .C(n394), .Z(n525) );
  GTECH_NAND2 U574 ( .A(n12), .B(n400), .Z(n394) );
  GTECH_NOT U575 ( .A(n11), .Z(n286) );
  GTECH_NOT U576 ( .A(n266), .Z(n524) );
  GTECH_NOT U577 ( .A(n295), .Z(n287) );
  GTECH_NAND2 U578 ( .A(N82), .B(n10), .Z(n295) );
  GTECH_NOT U579 ( .A(n526), .Z(N82) );
  GTECH_NOT U580 ( .A(n29), .Z(n388) );
  GTECH_NOT U581 ( .A(n527), .Z(n285) );
  GTECH_MUX2 U582 ( .A(n526), .B(n528), .S(n10), .Z(n527) );
  GTECH_NAND2 U583 ( .A(n28), .B(n296), .Z(n528) );
  GTECH_NAND2 U584 ( .A(n296), .B(n404), .Z(n526) );
  GTECH_NOT U585 ( .A(n28), .Z(n404) );
  GTECH_NOT U586 ( .A(n294), .Z(n283) );
  GTECH_NAND3 U587 ( .A(n296), .B(n402), .C(n28), .Z(n294) );
  GTECH_NOT U588 ( .A(n10), .Z(n402) );
  GTECH_NOT U589 ( .A(n318), .Z(n296) );
  GTECH_OAI21 U590 ( .A(n314), .B(n315), .C(n529), .Z(n318) );
  GTECH_AND2 U591 ( .A(n316), .B(n317), .Z(n529) );
  GTECH_NOT U592 ( .A(Rst), .Z(n317) );
  GTECH_NOT U593 ( .A(Ld), .Z(n316) );
  GTECH_NOT U594 ( .A(n9), .Z(n315) );
  GTECH_NAND2 U595 ( .A(n8), .B(n320), .Z(n314) );
  GTECH_NOT U596 ( .A(n323), .Z(n320) );
  GTECH_NAND2 U597 ( .A(n7), .B(n322), .Z(n323) );
  GTECH_NOT U598 ( .A(n530), .Z(n322) );
  GTECH_NAND2 U599 ( .A(n6), .B(n264), .Z(n530) );
  GTECH_XOR2 U600 ( .A(n522), .B(n514), .Z(n387) );
  GTECH_ADD_ABC U601 ( .A(n266), .B(n11), .C(n398), .COUT(n514) );
  GTECH_NAND2 U602 ( .A(n290), .B(n400), .Z(n398) );
  GTECH_NOT U603 ( .A(n265), .Z(n400) );
  GTECH_NOT U604 ( .A(n12), .Z(n290) );
  GTECH_XOR2 U605 ( .A(n517), .B(n29), .Z(n522) );
  GTECH_NOT U606 ( .A(n267), .Z(n517) );
endmodule

